LIBRARY IEEE; 
  USE IEEE.std_logic_1164.all; 
  USE IEEE.numeric_std.all; 

ENTITY COREDDS_C0_COREDDS_C0_0_dds_qrtr_cos IS 
  PORT ( 
    index : IN std_logic_vector(8 DOWNTO 0); 
    cosine : OUT std_logic_vector(11 DOWNTO 0)); 

    attribute syn_noclockbuf: Boolean;                     
    attribute syn_noclockbuf of index   : signal is true;  
    attribute syn_noclockbuf of cosine  : signal is true;  
END ENTITY COREDDS_C0_COREDDS_C0_0_dds_qrtr_cos; 

ARCHITECTURE rtl OF COREDDS_C0_COREDDS_C0_0_dds_qrtr_cos IS 
  SIGNAL A_int : integer; 
BEGIN 
  A_int <= to_integer(unsigned(index)); 
  PROCESS (A_int) 
    VARIABLE wave : std_logic_vector(11 DOWNTO 0); 
  BEGIN 
    CASE A_int IS      -- synopsys parallel_case     
      WHEN    0 => wave := "010000000000"; --        724 
      WHEN    1 => wave := "010000000000"; --        724 
      WHEN    2 => wave := "010000000000"; --        724 
      WHEN    3 => wave := "010000000000"; --        724 
      WHEN    4 => wave := "010000000000"; --        724 
      WHEN    5 => wave := "010000000000"; --        724 
      WHEN    6 => wave := "010000000000"; --        724 
      WHEN    7 => wave := "010000000000"; --        724 
      WHEN    8 => wave := "010000000000"; --        724 
      WHEN    9 => wave := "010000000000"; --        724 
      WHEN   10 => wave := "010000000000"; --        724 
      WHEN   11 => wave := "010000000000"; --        724 
      WHEN   12 => wave := "010000000000"; --        724 
      WHEN   13 => wave := "010000000000"; --        724 
      WHEN   14 => wave := "010000000000"; --        724 
      WHEN   15 => wave := "010000000000"; --        724 
      WHEN   16 => wave := "010000000000"; --        724 
      WHEN   17 => wave := "010000000000"; --        724 
      WHEN   18 => wave := "010000000000"; --        724 
      WHEN   19 => wave := "010000000000"; --        724 
      WHEN   20 => wave := "001111111111"; --        724 
      WHEN   21 => wave := "001111111111"; --        724 
      WHEN   22 => wave := "001111111111"; --        724 
      WHEN   23 => wave := "001111111111"; --        724 
      WHEN   24 => wave := "001111111111"; --        724 
      WHEN   25 => wave := "001111111111"; --        724 
      WHEN   26 => wave := "001111111111"; --        724 
      WHEN   27 => wave := "001111111111"; --        724 
      WHEN   28 => wave := "001111111111"; --        724 
      WHEN   29 => wave := "001111111111"; --        724 
      WHEN   30 => wave := "001111111111"; --        724 
      WHEN   31 => wave := "001111111111"; --        724 
      WHEN   32 => wave := "001111111111"; --        724 
      WHEN   33 => wave := "001111111111"; --        724 
      WHEN   34 => wave := "001111111111"; --        724 
      WHEN   35 => wave := "001111111110"; --        724 
      WHEN   36 => wave := "001111111110"; --        724 
      WHEN   37 => wave := "001111111110"; --        724 
      WHEN   38 => wave := "001111111110"; --        724 
      WHEN   39 => wave := "001111111110"; --        724 
      WHEN   40 => wave := "001111111110"; --        724 
      WHEN   41 => wave := "001111111110"; --        724 
      WHEN   42 => wave := "001111111110"; --        724 
      WHEN   43 => wave := "001111111110"; --        724 
      WHEN   44 => wave := "001111111110"; --        724 
      WHEN   45 => wave := "001111111110"; --        724 
      WHEN   46 => wave := "001111111101"; --        724 
      WHEN   47 => wave := "001111111101"; --        724 
      WHEN   48 => wave := "001111111101"; --        724 
      WHEN   49 => wave := "001111111101"; --        724 
      WHEN   50 => wave := "001111111101"; --        724 
      WHEN   51 => wave := "001111111101"; --        724 
      WHEN   52 => wave := "001111111101"; --        724 
      WHEN   53 => wave := "001111111101"; --        724 
      WHEN   54 => wave := "001111111100"; --        724 
      WHEN   55 => wave := "001111111100"; --        724 
      WHEN   56 => wave := "001111111100"; --        724 
      WHEN   57 => wave := "001111111100"; --        724 
      WHEN   58 => wave := "001111111100"; --        724 
      WHEN   59 => wave := "001111111100"; --        724 
      WHEN   60 => wave := "001111111100"; --        724 
      WHEN   61 => wave := "001111111011"; --        724 
      WHEN   62 => wave := "001111111011"; --        724 
      WHEN   63 => wave := "001111111011"; --        724 
      WHEN   64 => wave := "001111111011"; --        724 
      WHEN   65 => wave := "001111111011"; --        724 
      WHEN   66 => wave := "001111111011"; --        724 
      WHEN   67 => wave := "001111111011"; --        724 
      WHEN   68 => wave := "001111111010"; --        724 
      WHEN   69 => wave := "001111111010"; --        724 
      WHEN   70 => wave := "001111111010"; --        724 
      WHEN   71 => wave := "001111111010"; --        724 
      WHEN   72 => wave := "001111111010"; --        724 
      WHEN   73 => wave := "001111111001"; --        724 
      WHEN   74 => wave := "001111111001"; --        724 
      WHEN   75 => wave := "001111111001"; --        724 
      WHEN   76 => wave := "001111111001"; --        724 
      WHEN   77 => wave := "001111111001"; --        724 
      WHEN   78 => wave := "001111111001"; --        724 
      WHEN   79 => wave := "001111111000"; --        724 
      WHEN   80 => wave := "001111111000"; --        724 
      WHEN   81 => wave := "001111111000"; --        724 
      WHEN   82 => wave := "001111111000"; --        724 
      WHEN   83 => wave := "001111111000"; --        724 
      WHEN   84 => wave := "001111110111"; --        724 
      WHEN   85 => wave := "001111110111"; --        724 
      WHEN   86 => wave := "001111110111"; --        724 
      WHEN   87 => wave := "001111110111"; --        724 
      WHEN   88 => wave := "001111110111"; --        724 
      WHEN   89 => wave := "001111110110"; --        724 
      WHEN   90 => wave := "001111110110"; --        724 
      WHEN   91 => wave := "001111110110"; --        724 
      WHEN   92 => wave := "001111110110"; --        724 
      WHEN   93 => wave := "001111110101"; --        724 
      WHEN   94 => wave := "001111110101"; --        724 
      WHEN   95 => wave := "001111110101"; --        724 
      WHEN   96 => wave := "001111110101"; --        724 
      WHEN   97 => wave := "001111110101"; --        724 
      WHEN   98 => wave := "001111110100"; --        724 
      WHEN   99 => wave := "001111110100"; --        724 
      WHEN  100 => wave := "001111110100"; --        724 
      WHEN  101 => wave := "001111110100"; --        724 
      WHEN  102 => wave := "001111110011"; --        724 
      WHEN  103 => wave := "001111110011"; --        724 
      WHEN  104 => wave := "001111110011"; --        724 
      WHEN  105 => wave := "001111110011"; --        724 
      WHEN  106 => wave := "001111110010"; --        724 
      WHEN  107 => wave := "001111110010"; --        724 
      WHEN  108 => wave := "001111110010"; --        724 
      WHEN  109 => wave := "001111110010"; --        724 
      WHEN  110 => wave := "001111110001"; --        724 
      WHEN  111 => wave := "001111110001"; --        724 
      WHEN  112 => wave := "001111110001"; --        724 
      WHEN  113 => wave := "001111110001"; --        724 
      WHEN  114 => wave := "001111110000"; --        724 
      WHEN  115 => wave := "001111110000"; --        724 
      WHEN  116 => wave := "001111110000"; --        724 
      WHEN  117 => wave := "001111101111"; --        724 
      WHEN  118 => wave := "001111101111"; --        724 
      WHEN  119 => wave := "001111101111"; --        724 
      WHEN  120 => wave := "001111101111"; --        724 
      WHEN  121 => wave := "001111101110"; --        724 
      WHEN  122 => wave := "001111101110"; --        724 
      WHEN  123 => wave := "001111101110"; --        724 
      WHEN  124 => wave := "001111101101"; --        724 
      WHEN  125 => wave := "001111101101"; --        724 
      WHEN  126 => wave := "001111101101"; --        724 
      WHEN  127 => wave := "001111101100"; --        724 
      WHEN  128 => wave := "001111101100"; --        724 
      WHEN  129 => wave := "001111101100"; --        724 
      WHEN  130 => wave := "001111101100"; --        724 
      WHEN  131 => wave := "001111101011"; --        724 
      WHEN  132 => wave := "001111101011"; --        724 
      WHEN  133 => wave := "001111101011"; --        724 
      WHEN  134 => wave := "001111101010"; --        724 
      WHEN  135 => wave := "001111101010"; --        724 
      WHEN  136 => wave := "001111101010"; --        724 
      WHEN  137 => wave := "001111101001"; --        724 
      WHEN  138 => wave := "001111101001"; --        724 
      WHEN  139 => wave := "001111101001"; --        724 
      WHEN  140 => wave := "001111101000"; --        724 
      WHEN  141 => wave := "001111101000"; --        724 
      WHEN  142 => wave := "001111101000"; --        724 
      WHEN  143 => wave := "001111100111"; --        724 
      WHEN  144 => wave := "001111100111"; --        724 
      WHEN  145 => wave := "001111100111"; --        724 
      WHEN  146 => wave := "001111100110"; --        724 
      WHEN  147 => wave := "001111100110"; --        724 
      WHEN  148 => wave := "001111100110"; --        724 
      WHEN  149 => wave := "001111100101"; --        724 
      WHEN  150 => wave := "001111100101"; --        724 
      WHEN  151 => wave := "001111100100"; --        724 
      WHEN  152 => wave := "001111100100"; --        724 
      WHEN  153 => wave := "001111100100"; --        724 
      WHEN  154 => wave := "001111100011"; --        724 
      WHEN  155 => wave := "001111100011"; --        724 
      WHEN  156 => wave := "001111100011"; --        724 
      WHEN  157 => wave := "001111100010"; --        724 
      WHEN  158 => wave := "001111100010"; --        724 
      WHEN  159 => wave := "001111100010"; --        724 
      WHEN  160 => wave := "001111100001"; --        724 
      WHEN  161 => wave := "001111100001"; --        724 
      WHEN  162 => wave := "001111100000"; --        724 
      WHEN  163 => wave := "001111100000"; --        724 
      WHEN  164 => wave := "001111100000"; --        724 
      WHEN  165 => wave := "001111011111"; --        724 
      WHEN  166 => wave := "001111011111"; --        724 
      WHEN  167 => wave := "001111011110"; --        724 
      WHEN  168 => wave := "001111011110"; --        724 
      WHEN  169 => wave := "001111011110"; --        724 
      WHEN  170 => wave := "001111011101"; --        724 
      WHEN  171 => wave := "001111011101"; --        724 
      WHEN  172 => wave := "001111011100"; --        724 
      WHEN  173 => wave := "001111011100"; --        724 
      WHEN  174 => wave := "001111011100"; --        724 
      WHEN  175 => wave := "001111011011"; --        724 
      WHEN  176 => wave := "001111011011"; --        724 
      WHEN  177 => wave := "001111011010"; --        724 
      WHEN  178 => wave := "001111011010"; --        724 
      WHEN  179 => wave := "001111011001"; --        724 
      WHEN  180 => wave := "001111011001"; --        724 
      WHEN  181 => wave := "001111011001"; --        724 
      WHEN  182 => wave := "001111011000"; --        724 
      WHEN  183 => wave := "001111011000"; --        724 
      WHEN  184 => wave := "001111010111"; --        724 
      WHEN  185 => wave := "001111010111"; --        724 
      WHEN  186 => wave := "001111010110"; --        724 
      WHEN  187 => wave := "001111010110"; --        724 
      WHEN  188 => wave := "001111010101"; --        724 
      WHEN  189 => wave := "001111010101"; --        724 
      WHEN  190 => wave := "001111010101"; --        724 
      WHEN  191 => wave := "001111010100"; --        724 
      WHEN  192 => wave := "001111010100"; --        724 
      WHEN  193 => wave := "001111010011"; --        724 
      WHEN  194 => wave := "001111010011"; --        724 
      WHEN  195 => wave := "001111010010"; --        724 
      WHEN  196 => wave := "001111010010"; --        724 
      WHEN  197 => wave := "001111010001"; --        724 
      WHEN  198 => wave := "001111010001"; --        724 
      WHEN  199 => wave := "001111010000"; --        724 
      WHEN  200 => wave := "001111010000"; --        724 
      WHEN  201 => wave := "001111001111"; --        724 
      WHEN  202 => wave := "001111001111"; --        724 
      WHEN  203 => wave := "001111001111"; --        724 
      WHEN  204 => wave := "001111001110"; --        724 
      WHEN  205 => wave := "001111001110"; --        724 
      WHEN  206 => wave := "001111001101"; --        724 
      WHEN  207 => wave := "001111001101"; --        724 
      WHEN  208 => wave := "001111001100"; --        724 
      WHEN  209 => wave := "001111001100"; --        724 
      WHEN  210 => wave := "001111001011"; --        724 
      WHEN  211 => wave := "001111001011"; --        724 
      WHEN  212 => wave := "001111001010"; --        724 
      WHEN  213 => wave := "001111001010"; --        724 
      WHEN  214 => wave := "001111001001"; --        724 
      WHEN  215 => wave := "001111001001"; --        724 
      WHEN  216 => wave := "001111001000"; --        724 
      WHEN  217 => wave := "001111001000"; --        724 
      WHEN  218 => wave := "001111000111"; --        724 
      WHEN  219 => wave := "001111000110"; --        724 
      WHEN  220 => wave := "001111000110"; --        724 
      WHEN  221 => wave := "001111000101"; --        724 
      WHEN  222 => wave := "001111000101"; --        724 
      WHEN  223 => wave := "001111000100"; --        724 
      WHEN  224 => wave := "001111000100"; --        724 
      WHEN  225 => wave := "001111000011"; --        724 
      WHEN  226 => wave := "001111000011"; --        724 
      WHEN  227 => wave := "001111000010"; --        724 
      WHEN  228 => wave := "001111000010"; --        724 
      WHEN  229 => wave := "001111000001"; --        724 
      WHEN  230 => wave := "001111000001"; --        724 
      WHEN  231 => wave := "001111000000"; --        724 
      WHEN  232 => wave := "001111000000"; --        724 
      WHEN  233 => wave := "001110111111"; --        724 
      WHEN  234 => wave := "001110111110"; --        724 
      WHEN  235 => wave := "001110111110"; --        724 
      WHEN  236 => wave := "001110111101"; --        724 
      WHEN  237 => wave := "001110111101"; --        724 
      WHEN  238 => wave := "001110111100"; --        724 
      WHEN  239 => wave := "001110111100"; --        724 
      WHEN  240 => wave := "001110111011"; --        724 
      WHEN  241 => wave := "001110111011"; --        724 
      WHEN  242 => wave := "001110111010"; --        724 
      WHEN  243 => wave := "001110111001"; --        724 
      WHEN  244 => wave := "001110111001"; --        724 
      WHEN  245 => wave := "001110111000"; --        724 
      WHEN  246 => wave := "001110111000"; --        724 
      WHEN  247 => wave := "001110110111"; --        724 
      WHEN  248 => wave := "001110110110"; --        724 
      WHEN  249 => wave := "001110110110"; --        724 
      WHEN  250 => wave := "001110110101"; --        724 
      WHEN  251 => wave := "001110110101"; --        724 
      WHEN  252 => wave := "001110110100"; --        724 
      WHEN  253 => wave := "001110110100"; --        724 
      WHEN  254 => wave := "001110110011"; --        724 
      WHEN  255 => wave := "001110110010"; --        724 
      WHEN  256 => wave := "001110110010"; --        724 
      WHEN  257 => wave := "001110110001"; --        724 
      WHEN  258 => wave := "001110110001"; --        724 
      WHEN  259 => wave := "001110110000"; --        724 
      WHEN  260 => wave := "001110101111"; --        724 
      WHEN  261 => wave := "001110101111"; --        724 
      WHEN  262 => wave := "001110101110"; --        724 
      WHEN  263 => wave := "001110101101"; --        724 
      WHEN  264 => wave := "001110101101"; --        724 
      WHEN  265 => wave := "001110101100"; --        724 
      WHEN  266 => wave := "001110101100"; --        724 
      WHEN  267 => wave := "001110101011"; --        724 
      WHEN  268 => wave := "001110101010"; --        724 
      WHEN  269 => wave := "001110101010"; --        724 
      WHEN  270 => wave := "001110101001"; --        724 
      WHEN  271 => wave := "001110101000"; --        724 
      WHEN  272 => wave := "001110101000"; --        724 
      WHEN  273 => wave := "001110100111"; --        724 
      WHEN  274 => wave := "001110100111"; --        724 
      WHEN  275 => wave := "001110100110"; --        724 
      WHEN  276 => wave := "001110100101"; --        724 
      WHEN  277 => wave := "001110100101"; --        724 
      WHEN  278 => wave := "001110100100"; --        724 
      WHEN  279 => wave := "001110100011"; --        724 
      WHEN  280 => wave := "001110100011"; --        724 
      WHEN  281 => wave := "001110100010"; --        724 
      WHEN  282 => wave := "001110100001"; --        724 
      WHEN  283 => wave := "001110100001"; --        724 
      WHEN  284 => wave := "001110100000"; --        724 
      WHEN  285 => wave := "001110011111"; --        724 
      WHEN  286 => wave := "001110011111"; --        724 
      WHEN  287 => wave := "001110011110"; --        724 
      WHEN  288 => wave := "001110011101"; --        724 
      WHEN  289 => wave := "001110011101"; --        724 
      WHEN  290 => wave := "001110011100"; --        724 
      WHEN  291 => wave := "001110011011"; --        724 
      WHEN  292 => wave := "001110011011"; --        724 
      WHEN  293 => wave := "001110011010"; --        724 
      WHEN  294 => wave := "001110011001"; --        724 
      WHEN  295 => wave := "001110011001"; --        724 
      WHEN  296 => wave := "001110011000"; --        724 
      WHEN  297 => wave := "001110010111"; --        724 
      WHEN  298 => wave := "001110010111"; --        724 
      WHEN  299 => wave := "001110010110"; --        724 
      WHEN  300 => wave := "001110010101"; --        724 
      WHEN  301 => wave := "001110010100"; --        724 
      WHEN  302 => wave := "001110010100"; --        724 
      WHEN  303 => wave := "001110010011"; --        724 
      WHEN  304 => wave := "001110010010"; --        724 
      WHEN  305 => wave := "001110010010"; --        724 
      WHEN  306 => wave := "001110010001"; --        724 
      WHEN  307 => wave := "001110010000"; --        724 
      WHEN  308 => wave := "001110001111"; --        724 
      WHEN  309 => wave := "001110001111"; --        724 
      WHEN  310 => wave := "001110001110"; --        724 
      WHEN  311 => wave := "001110001101"; --        724 
      WHEN  312 => wave := "001110001101"; --        724 
      WHEN  313 => wave := "001110001100"; --        724 
      WHEN  314 => wave := "001110001011"; --        724 
      WHEN  315 => wave := "001110001010"; --        724 
      WHEN  316 => wave := "001110001010"; --        724 
      WHEN  317 => wave := "001110001001"; --        724 
      WHEN  318 => wave := "001110001000"; --        724 
      WHEN  319 => wave := "001110000111"; --        724 
      WHEN  320 => wave := "001110000111"; --        724 
      WHEN  321 => wave := "001110000110"; --        724 
      WHEN  322 => wave := "001110000101"; --        724 
      WHEN  323 => wave := "001110000100"; --        724 
      WHEN  324 => wave := "001110000100"; --        724 
      WHEN  325 => wave := "001110000011"; --        724 
      WHEN  326 => wave := "001110000010"; --        724 
      WHEN  327 => wave := "001110000001"; --        724 
      WHEN  328 => wave := "001110000001"; --        724 
      WHEN  329 => wave := "001110000000"; --        724 
      WHEN  330 => wave := "001101111111"; --        724 
      WHEN  331 => wave := "001101111110"; --        724 
      WHEN  332 => wave := "001101111110"; --        724 
      WHEN  333 => wave := "001101111101"; --        724 
      WHEN  334 => wave := "001101111100"; --        724 
      WHEN  335 => wave := "001101111011"; --        724 
      WHEN  336 => wave := "001101111011"; --        724 
      WHEN  337 => wave := "001101111010"; --        724 
      WHEN  338 => wave := "001101111001"; --        724 
      WHEN  339 => wave := "001101111000"; --        724 
      WHEN  340 => wave := "001101110111"; --        724 
      WHEN  341 => wave := "001101110111"; --        724 
      WHEN  342 => wave := "001101110110"; --        724 
      WHEN  343 => wave := "001101110101"; --        724 
      WHEN  344 => wave := "001101110100"; --        724 
      WHEN  345 => wave := "001101110100"; --        724 
      WHEN  346 => wave := "001101110011"; --        724 
      WHEN  347 => wave := "001101110010"; --        724 
      WHEN  348 => wave := "001101110001"; --        724 
      WHEN  349 => wave := "001101110000"; --        724 
      WHEN  350 => wave := "001101110000"; --        724 
      WHEN  351 => wave := "001101101111"; --        724 
      WHEN  352 => wave := "001101101110"; --        724 
      WHEN  353 => wave := "001101101101"; --        724 
      WHEN  354 => wave := "001101101100"; --        724 
      WHEN  355 => wave := "001101101011"; --        724 
      WHEN  356 => wave := "001101101011"; --        724 
      WHEN  357 => wave := "001101101010"; --        724 
      WHEN  358 => wave := "001101101001"; --        724 
      WHEN  359 => wave := "001101101000"; --        724 
      WHEN  360 => wave := "001101100111"; --        724 
      WHEN  361 => wave := "001101100111"; --        724 
      WHEN  362 => wave := "001101100110"; --        724 
      WHEN  363 => wave := "001101100101"; --        724 
      WHEN  364 => wave := "001101100100"; --        724 
      WHEN  365 => wave := "001101100011"; --        724 
      WHEN  366 => wave := "001101100010"; --        724 
      WHEN  367 => wave := "001101100010"; --        724 
      WHEN  368 => wave := "001101100001"; --        724 
      WHEN  369 => wave := "001101100000"; --        724 
      WHEN  370 => wave := "001101011111"; --        724 
      WHEN  371 => wave := "001101011110"; --        724 
      WHEN  372 => wave := "001101011101"; --        724 
      WHEN  373 => wave := "001101011100"; --        724 
      WHEN  374 => wave := "001101011100"; --        724 
      WHEN  375 => wave := "001101011011"; --        724 
      WHEN  376 => wave := "001101011010"; --        724 
      WHEN  377 => wave := "001101011001"; --        724 
      WHEN  378 => wave := "001101011000"; --        724 
      WHEN  379 => wave := "001101010111"; --        724 
      WHEN  380 => wave := "001101010110"; --        724 
      WHEN  381 => wave := "001101010110"; --        724 
      WHEN  382 => wave := "001101010101"; --        724 
      WHEN  383 => wave := "001101010100"; --        724 
      WHEN  384 => wave := "001101010011"; --        724 
      WHEN  385 => wave := "001101010010"; --        724 
      WHEN  386 => wave := "001101010001"; --        724 
      WHEN  387 => wave := "001101010000"; --        724 
      WHEN  388 => wave := "001101001111"; --        724 
      WHEN  389 => wave := "001101001111"; --        724 
      WHEN  390 => wave := "001101001110"; --        724 
      WHEN  391 => wave := "001101001101"; --        724 
      WHEN  392 => wave := "001101001100"; --        724 
      WHEN  393 => wave := "001101001011"; --        724 
      WHEN  394 => wave := "001101001010"; --        724 
      WHEN  395 => wave := "001101001001"; --        724 
      WHEN  396 => wave := "001101001000"; --        724 
      WHEN  397 => wave := "001101000111"; --        724 
      WHEN  398 => wave := "001101000111"; --        724 
      WHEN  399 => wave := "001101000110"; --        724 
      WHEN  400 => wave := "001101000101"; --        724 
      WHEN  401 => wave := "001101000100"; --        724 
      WHEN  402 => wave := "001101000011"; --        724 
      WHEN  403 => wave := "001101000010"; --        724 
      WHEN  404 => wave := "001101000001"; --        724 
      WHEN  405 => wave := "001101000000"; --        724 
      WHEN  406 => wave := "001100111111"; --        724 
      WHEN  407 => wave := "001100111110"; --        724 
      WHEN  408 => wave := "001100111101"; --        724 
      WHEN  409 => wave := "001100111101"; --        724 
      WHEN  410 => wave := "001100111100"; --        724 
      WHEN  411 => wave := "001100111011"; --        724 
      WHEN  412 => wave := "001100111010"; --        724 
      WHEN  413 => wave := "001100111001"; --        724 
      WHEN  414 => wave := "001100111000"; --        724 
      WHEN  415 => wave := "001100110111"; --        724 
      WHEN  416 => wave := "001100110110"; --        724 
      WHEN  417 => wave := "001100110101"; --        724 
      WHEN  418 => wave := "001100110100"; --        724 
      WHEN  419 => wave := "001100110011"; --        724 
      WHEN  420 => wave := "001100110010"; --        724 
      WHEN  421 => wave := "001100110001"; --        724 
      WHEN  422 => wave := "001100110000"; --        724 
      WHEN  423 => wave := "001100101111"; --        724 
      WHEN  424 => wave := "001100101110"; --        724 
      WHEN  425 => wave := "001100101110"; --        724 
      WHEN  426 => wave := "001100101101"; --        724 
      WHEN  427 => wave := "001100101100"; --        724 
      WHEN  428 => wave := "001100101011"; --        724 
      WHEN  429 => wave := "001100101010"; --        724 
      WHEN  430 => wave := "001100101001"; --        724 
      WHEN  431 => wave := "001100101000"; --        724 
      WHEN  432 => wave := "001100100111"; --        724 
      WHEN  433 => wave := "001100100110"; --        724 
      WHEN  434 => wave := "001100100101"; --        724 
      WHEN  435 => wave := "001100100100"; --        724 
      WHEN  436 => wave := "001100100011"; --        724 
      WHEN  437 => wave := "001100100010"; --        724 
      WHEN  438 => wave := "001100100001"; --        724 
      WHEN  439 => wave := "001100100000"; --        724 
      WHEN  440 => wave := "001100011111"; --        724 
      WHEN  441 => wave := "001100011110"; --        724 
      WHEN  442 => wave := "001100011101"; --        724 
      WHEN  443 => wave := "001100011100"; --        724 
      WHEN  444 => wave := "001100011011"; --        724 
      WHEN  445 => wave := "001100011010"; --        724 
      WHEN  446 => wave := "001100011001"; --        724 
      WHEN  447 => wave := "001100011000"; --        724 
      WHEN  448 => wave := "001100010111"; --        724 
      WHEN  449 => wave := "001100010110"; --        724 
      WHEN  450 => wave := "001100010101"; --        724 
      WHEN  451 => wave := "001100010100"; --        724 
      WHEN  452 => wave := "001100010011"; --        724 
      WHEN  453 => wave := "001100010010"; --        724 
      WHEN  454 => wave := "001100010001"; --        724 
      WHEN  455 => wave := "001100010000"; --        724 
      WHEN  456 => wave := "001100001111"; --        724 
      WHEN  457 => wave := "001100001110"; --        724 
      WHEN  458 => wave := "001100001101"; --        724 
      WHEN  459 => wave := "001100001100"; --        724 
      WHEN  460 => wave := "001100001011"; --        724 
      WHEN  461 => wave := "001100001010"; --        724 
      WHEN  462 => wave := "001100001001"; --        724 
      WHEN  463 => wave := "001100001000"; --        724 
      WHEN  464 => wave := "001100000111"; --        724 
      WHEN  465 => wave := "001100000110"; --        724 
      WHEN  466 => wave := "001100000101"; --        724 
      WHEN  467 => wave := "001100000100"; --        724 
      WHEN  468 => wave := "001100000011"; --        724 
      WHEN  469 => wave := "001100000010"; --        724 
      WHEN  470 => wave := "001100000001"; --        724 
      WHEN  471 => wave := "001100000000"; --        724 
      WHEN  472 => wave := "001011111111"; --        724 
      WHEN  473 => wave := "001011111110"; --        724 
      WHEN  474 => wave := "001011111101"; --        724 
      WHEN  475 => wave := "001011111011"; --        724 
      WHEN  476 => wave := "001011111010"; --        724 
      WHEN  477 => wave := "001011111001"; --        724 
      WHEN  478 => wave := "001011111000"; --        724 
      WHEN  479 => wave := "001011110111"; --        724 
      WHEN  480 => wave := "001011110110"; --        724 
      WHEN  481 => wave := "001011110101"; --        724 
      WHEN  482 => wave := "001011110100"; --        724 
      WHEN  483 => wave := "001011110011"; --        724 
      WHEN  484 => wave := "001011110010"; --        724 
      WHEN  485 => wave := "001011110001"; --        724 
      WHEN  486 => wave := "001011110000"; --        724 
      WHEN  487 => wave := "001011101111"; --        724 
      WHEN  488 => wave := "001011101110"; --        724 
      WHEN  489 => wave := "001011101101"; --        724 
      WHEN  490 => wave := "001011101100"; --        724 
      WHEN  491 => wave := "001011101010"; --        724 
      WHEN  492 => wave := "001011101001"; --        724 
      WHEN  493 => wave := "001011101000"; --        724 
      WHEN  494 => wave := "001011100111"; --        724 
      WHEN  495 => wave := "001011100110"; --        724 
      WHEN  496 => wave := "001011100101"; --        724 
      WHEN  497 => wave := "001011100100"; --        724 
      WHEN  498 => wave := "001011100011"; --        724 
      WHEN  499 => wave := "001011100010"; --        724 
      WHEN  500 => wave := "001011100001"; --        724 
      WHEN  501 => wave := "001011100000"; --        724 
      WHEN  502 => wave := "001011011111"; --        724 
      WHEN  503 => wave := "001011011101"; --        724 
      WHEN  504 => wave := "001011011100"; --        724 
      WHEN  505 => wave := "001011011011"; --        724 
      WHEN  506 => wave := "001011011010"; --        724 
      WHEN  507 => wave := "001011011001"; --        724 
      WHEN  508 => wave := "001011011000"; --        724 
      WHEN  509 => wave := "001011010111"; --        724 
      WHEN  510 => wave := "001011010110"; --        724 
      WHEN OTHERS => wave := "001011010101"; --        725 
    END CASE; 

    cosine <= wave; 

  END PROCESS; 
END ARCHITECTURE rtl; 
