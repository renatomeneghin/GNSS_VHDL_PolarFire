-- -----------------------------------------------------------------------------
--Actel Corporation Proprietary and Confidential
--Copyright 2008 Actel Corporation. All rights reserved.
--
--ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
--ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
--IN ADVANCE IN WRITING.
--
--Description:  CoreFFT Test bench 
--              Input/Output golden test vectors 
--
--Revision Information:
--Date         Description
--05Nov2009    Initial Release 
--
--SVN Revision Information:
--SVN $Revision: $
--SVN $Data: $
--
--Resolved SARs
--SAR     Date    Who         Description
--
--Notes:

-----------------------------------------------------------
LIBRARY IEEE; 
  USE IEEE.std_logic_1164.all; 

ENTITY testvect1 IS 
  PORT ( 
    A : IN integer; 
    T : OUT std_logic_vector(47 DOWNTO 0));
END ENTITY testvect1; 

ARCHITECTURE arch_rom OF testvect1 IS 
BEGIN 
  PROCESS (A) 
    VARIABLE Ti  : std_logic_vector(47 DOWNTO 0); 
  BEGIN 
    CASE A IS  
      WHEN    0 => Ti := "000000000000000000000000011001100110011001100101"; --         +0   +6710885
      WHEN    1 => Ti := "000000001010000011011001011001100110010111100111"; --     +41177   +6710759
      WHEN    2 => Ti := "000000010100000110110000011001100110010001101100"; --     +82352   +6710380
      WHEN    3 => Ti := "000000011110001010000101011001100110000111110100"; --    +123525   +6709748
      WHEN    4 => Ti := "000000101000001101010101011001100101111010000000"; --    +164693   +6708864
      WHEN    5 => Ti := "000000110010010000011111011001100101101000001111"; --    +205855   +6707727
      WHEN    6 => Ti := "000000111100010011100001011001100101010010100010"; --    +247009   +6706338
      WHEN    7 => Ti := "000001000110010110011001011001100100111000111000"; --    +288153   +6704696
      WHEN    8 => Ti := "000001010000011001000111011001100100011011010010"; --    +329287   +6702802
      WHEN    9 => Ti := "000001011010011011101000011001100011111001101111"; --    +370408   +6700655
      WHEN   10 => Ti := "000001100100011101111100011001100011010100010000"; --    +411516   +6698256
      WHEN   11 => Ti := "000001101110100000000000011001100010101010110101"; --    +452608   +6695605
      WHEN   12 => Ti := "000001111000100001110011011001100001111101011110"; --    +493683   +6692702
      WHEN   13 => Ti := "000010000010100011010011011001100001001100001010"; --    +534739   +6689546
      WHEN   14 => Ti := "000010001100100100011111011001100000010110111011"; --    +575775   +6686139
      WHEN   15 => Ti := "000010010110100101010110011001011111011101110001"; --    +616790   +6682481
      WHEN   16 => Ti := "000010100000100101110101011001011110100000101010"; --    +657781   +6678570
      WHEN   17 => Ti := "000010101010100101111100011001011101011111101001"; --    +698748   +6674409
      WHEN   18 => Ti := "000010110100100101101000011001011100011010101011"; --    +739688   +6669995
      WHEN   19 => Ti := "000010111110100100111001011001011011010001110011"; --    +780601   +6665331
      WHEN   20 => Ti := "000011001000100011101100011001011010000101000000"; --    +821484   +6660416
      WHEN   21 => Ti := "000011010010100010000000011001011000110100010010"; --    +862336   +6655250
      WHEN   22 => Ti := "000011011100011111110011011001010111011111101010"; --    +903155   +6649834
      WHEN   23 => Ti := "000011100110011101000101011001010110000111000111"; --    +943941   +6644167
      WHEN   24 => Ti := "000011110000011001110011011001010100101010101010"; --    +984691   +6638250
      WHEN   25 => Ti := "000011111010010101111100011001010011001010010011"; --   +1025404   +6632083
      WHEN   26 => Ti := "000100000100010001011110011001010001100110000010"; --   +1066078   +6625666
      WHEN   27 => Ti := "000100001110001100011001011001001111111101111000"; --   +1106713   +6619000
      WHEN   28 => Ti := "000100011000000110101001011001001110010001110101"; --   +1147305   +6612085
      WHEN   29 => Ti := "000100100010000000001111011001001100100001111001"; --   +1187855   +6604921
      WHEN   30 => Ti := "000100101011111001000111011001001010101110000100"; --   +1228359   +6597508
      WHEN   31 => Ti := "000100110101110001010010011001001000110110010111"; --   +1268818   +6589847
      WHEN   32 => Ti := "000100111111101000101100011001000110111010110001"; --   +1309228   +6581937
      WHEN   33 => Ti := "000101001001011111010110011001000100111011010100"; --   +1349590   +6573780
      WHEN   34 => Ti := "000101010011010101001100011001000010110111111111"; --   +1389900   +6565375
      WHEN   35 => Ti := "000101011101001010001110011001000000110000110100"; --   +1430158   +6556724
      WHEN   36 => Ti := "000101100110111110011011011000111110100101110001"; --   +1470363   +6547825
      WHEN   37 => Ti := "000101110000110001110000011000111100010110111000"; --   +1510512   +6538680
      WHEN   38 => Ti := "000101111010100100001100011000111010000100001000"; --   +1550604   +6529288
      WHEN   39 => Ti := "000110000100010101101110011000110111101101100011"; --   +1590638   +6519651
      WHEN   40 => Ti := "000110001110000110010100011000110101010011001000"; --   +1630612   +6509768
      WHEN   41 => Ti := "000110010111110101111100011000110010110100111000"; --   +1670524   +6499640
      WHEN   42 => Ti := "000110100001100100100110011000110000010010110100"; --   +1710374   +6489268
      WHEN   43 => Ti := "000110101011010010001111011000101101101100111011"; --   +1750159   +6478651
      WHEN   44 => Ti := "000110110100111110110110011000101011000011001110"; --   +1789878   +6467790
      WHEN   45 => Ti := "000110111110101010011010011000101000010101101110"; --   +1829530   +6456686
      WHEN   46 => Ti := "000111001000010100111001011000100101100100011011"; --   +1869113   +6445339
      WHEN   47 => Ti := "000111010001111110010010011000100010101111010101"; --   +1908626   +6433749
      WHEN   48 => Ti := "000111011011100110100011011000011111110110011101"; --   +1948067   +6421917
      WHEN   49 => Ti := "000111100101001101101010011000011100111001110011"; --   +1987434   +6409843
      WHEN   50 => Ti := "000111101110110011100111011000011001111001010111"; --   +2026727   +6397527
      WHEN   51 => Ti := "000111111000011000010111011000010110110101001011"; --   +2065943   +6384971
      WHEN   52 => Ti := "001000000001111011111010011000010011101101001110"; --   +2105082   +6372174
      WHEN   53 => Ti := "001000001011011110001101011000010000100001100010"; --   +2144141   +6359138
      WHEN   54 => Ti := "001000010100111111010000011000001101010010000110"; --   +2183120   +6345862
      WHEN   55 => Ti := "001000011110011111000000011000001001111110111011"; --   +2222016   +6332347
      WHEN   56 => Ti := "001000100111111101011101011000000110101000000010"; --   +2260829   +6318594
      WHEN   57 => Ti := "001000110001011010100100011000000011001101011011"; --   +2299556   +6304603
      WHEN   58 => Ti := "001000111010110110010101010111111111101111000110"; --   +2338197   +6290374
      WHEN   59 => Ti := "001001000100010000101110010111111100001101000101"; --   +2376750   +6275909
      WHEN   60 => Ti := "001001001101101001101110010111111000100111010111"; --   +2415214   +6261207
      WHEN   61 => Ti := "001001010111000001010011010111110100111101111110"; --   +2453587   +6246270
      WHEN   62 => Ti := "001001100000010111011011010111110001010000111010"; --   +2491867   +6231098
      WHEN   63 => Ti := "001001101001101100000101010111101101100000001010"; --   +2530053   +6215690
      WHEN   64 => Ti := "001001110010111111010000010111101001101011110001"; --   +2568144   +6200049
      WHEN   65 => Ti := "001001111100010000111011010111100101110011101111"; --   +2606139   +6184175
      WHEN   66 => Ti := "001010000101100001000011010111100001111000000011"; --   +2644035   +6168067
      WHEN   67 => Ti := "001010001110101111101000010111011101111000110000"; --   +2681832   +6151728
      WHEN   68 => Ti := "001010010111111100101000010111011001110101110101"; --   +2719528   +6135157
      WHEN   69 => Ti := "001010100001001000000001010111010101101111010010"; --   +2757121   +6118354
      WHEN   70 => Ti := "001010101010010001110011010111010001100101001010"; --   +2794611   +6101322
      WHEN   71 => Ti := "001010110011011001111011010111001101010111011100"; --   +2831995   +6084060
      WHEN   72 => Ti := "001010111100100000011001010111001001000110001000"; --   +2869273   +6066568
      WHEN   73 => Ti := "001011000101100101001011010111000100110001010000"; --   +2906443   +6048848
      WHEN   74 => Ti := "001011001110101000001111010111000000011000110101"; --   +2943503   +6030901
      WHEN   75 => Ti := "001011010111101001100100010110111011111100110111"; --   +2980452   +6012727
      WHEN   76 => Ti := "001011100000101001001010010110110111011101010110"; --   +3017290   +5994326
      WHEN   77 => Ti := "001011101001100110111101010110110010111010010011"; --   +3054013   +5975699
      WHEN   78 => Ti := "001011110010100010111110010110101110010011101111"; --   +3090622   +5956847
      WHEN   79 => Ti := "001011111011011101001010010110101001101001101100"; --   +3127114   +5937772
      WHEN   80 => Ti := "001100000100010101100001010110100100111100001000"; --   +3163489   +5918472
      WHEN   81 => Ti := "001100001101001100000001010110100000001011000110"; --   +3199745   +5898950
      WHEN   82 => Ti := "001100010110000000101000010110011011010110100110"; --   +3235880   +5879206
      WHEN   83 => Ti := "001100011110110011010101010110010110011110101000"; --   +3271893   +5859240
      WHEN   84 => Ti := "001100100111100100000111010110010001100011001110"; --   +3307783   +5839054
      WHEN   85 => Ti := "001100110000010010111100010110001100100100011000"; --   +3343548   +5818648
      WHEN   86 => Ti := "001100111000111111110100010110000111100010000110"; --   +3379188   +5798022
      WHEN   87 => Ti := "001101000001101010101100010110000010011100011011"; --   +3414700   +5777179
      WHEN   88 => Ti := "001101001010010011100100010101111101010011010110"; --   +3450084   +5756118
      WHEN   89 => Ti := "001101010010111010011010010101111000000110111000"; --   +3485338   +5734840
      WHEN   90 => Ti := "001101011011011111001101010101110010110111000011"; --   +3520461   +5713347
      WHEN   91 => Ti := "001101100100000001111011010101101101100011110110"; --   +3555451   +5691638
      WHEN   92 => Ti := "001101101100100010100011010101101000001101010011"; --   +3590307   +5669715
      WHEN   93 => Ti := "001101110101000001000100010101100010110011011011"; --   +3625028   +5647579
      WHEN   94 => Ti := "001101111101011101011101010101011101010110001110"; --   +3659613   +5625230
      WHEN   95 => Ti := "001110000101110111101100010101010111110101101101"; --   +3694060   +5602669
      WHEN   96 => Ti := "001110001110001111110000010101010010010001111001"; --   +3728368   +5579897
      WHEN   97 => Ti := "001110010110100101100111010101001100101010110011"; --   +3762535   +5556915
      WHEN   98 => Ti := "001110011110111001010001010101000111000000011100"; --   +3796561   +5533724
      WHEN   99 => Ti := "001110100111001010101100010101000001010010110101"; --   +3830444   +5510325
      WHEN  100 => Ti := "001110101111011001110110010100111011100001111110"; --   +3864182   +5486718
      WHEN  101 => Ti := "001110110111100110110000010100110101101101111000"; --   +3897776   +5462904
      WHEN  102 => Ti := "001110111111110001010110010100101111110110100101"; --   +3931222   +5438885
      WHEN  103 => Ti := "001111000111111001101000010100101001111100000101"; --   +3964520   +5414661
      WHEN  104 => Ti := "001111001111111111100101010100100011111110011001"; --   +3997669   +5390233
      WHEN  105 => Ti := "001111011000000011001100010100011101111101100011"; --   +4030668   +5365603
      WHEN  106 => Ti := "001111100000000100011011010100010111111001100010"; --   +4063515   +5340770
      WHEN  107 => Ti := "001111101000000011010001010100010001110010011000"; --   +4096209   +5315736
      WHEN  108 => Ti := "001111101111111111101100010100001011101000000110"; --   +4128748   +5290502
      WHEN  109 => Ti := "001111110111111001101101010100000101011010101101"; --   +4161133   +5265069
      WHEN  110 => Ti := "001111111111110001010000010011111111001010001110"; --   +4193360   +5239438
      WHEN  111 => Ti := "010000000111100110010110010011111000110110101001"; --   +4225430   +5213609
      WHEN  112 => Ti := "010000001111011000111100010011110010100000000000"; --   +4257340   +5187584
      WHEN  113 => Ti := "010000010111001001000011010011101100000110010100"; --   +4289091   +5161364
      WHEN  114 => Ti := "010000011110110110100111010011100101101001100101"; --   +4320679   +5134949
      WHEN  115 => Ti := "010000100110100001101001010011011111001001110110"; --   +4352105   +5108342
      WHEN  116 => Ti := "010000101110001010001000010011011000100111000101"; --   +4383368   +5081541
      WHEN  117 => Ti := "010000110101110000000001010011010010000001010110"; --   +4414465   +5054550
      WHEN  118 => Ti := "010000111101010011010100010011001011011000101000"; --   +4445396   +5027368
      WHEN  119 => Ti := "010001000100110100000000010011000100101100111101"; --   +4476160   +4999997
      WHEN  120 => Ti := "010001001100010010000011010010111101111110010110"; --   +4506755   +4972438
      WHEN  121 => Ti := "010001010011101101011100010010110111001100110011"; --   +4537180   +4944691
      WHEN  122 => Ti := "010001011011000110001011010010110000011000010111"; --   +4567435   +4916759
      WHEN  123 => Ti := "010001100010011100001110010010101001100001000001"; --   +4597518   +4888641
      WHEN  124 => Ti := "010001101001101111100011010010100010100110110011"; --   +4627427   +4860339
      WHEN  125 => Ti := "010001110001000000001011010010011011101001101110"; --   +4657163   +4831854
      WHEN  126 => Ti := "010001111000001110000011010010010100101001110011"; --   +4686723   +4803187
      WHEN  127 => Ti := "010001111111011001001010010010001101100111000100"; --   +4716106   +4774340
      WHEN  128 => Ti := "010010000110100001100000010010000110100001100000"; --   +4745312   +4745312
      WHEN  129 => Ti := "010010001101100111000100010001111111011001001010"; --   +4774340   +4716106
      WHEN  130 => Ti := "010010010100101001110011010001111000001110000011"; --   +4803187   +4686723
      WHEN  131 => Ti := "010010011011101001101110010001110001000000001011"; --   +4831854   +4657163
      WHEN  132 => Ti := "010010100010100110110011010001101001101111100011"; --   +4860339   +4627427
      WHEN  133 => Ti := "010010101001100001000001010001100010011100001110"; --   +4888641   +4597518
      WHEN  134 => Ti := "010010110000011000010111010001011011000110001011"; --   +4916759   +4567435
      WHEN  135 => Ti := "010010110111001100110011010001010011101101011100"; --   +4944691   +4537180
      WHEN  136 => Ti := "010010111101111110010110010001001100010010000011"; --   +4972438   +4506755
      WHEN  137 => Ti := "010011000100101100111101010001000100110100000000"; --   +4999997   +4476160
      WHEN  138 => Ti := "010011001011011000101000010000111101010011010100"; --   +5027368   +4445396
      WHEN  139 => Ti := "010011010010000001010110010000110101110000000001"; --   +5054550   +4414465
      WHEN  140 => Ti := "010011011000100111000101010000101110001010001000"; --   +5081541   +4383368
      WHEN  141 => Ti := "010011011111001001110110010000100110100001101001"; --   +5108342   +4352105
      WHEN  142 => Ti := "010011100101101001100101010000011110110110100111"; --   +5134949   +4320679
      WHEN  143 => Ti := "010011101100000110010100010000010111001001000011"; --   +5161364   +4289091
      WHEN  144 => Ti := "010011110010100000000000010000001111011000111100"; --   +5187584   +4257340
      WHEN  145 => Ti := "010011111000110110101001010000000111100110010110"; --   +5213609   +4225430
      WHEN  146 => Ti := "010011111111001010001110001111111111110001010000"; --   +5239438   +4193360
      WHEN  147 => Ti := "010100000101011010101101001111110111111001101101"; --   +5265069   +4161133
      WHEN  148 => Ti := "010100001011101000000110001111101111111111101100"; --   +5290502   +4128748
      WHEN  149 => Ti := "010100010001110010011000001111101000000011010001"; --   +5315736   +4096209
      WHEN  150 => Ti := "010100010111111001100010001111100000000100011011"; --   +5340770   +4063515
      WHEN  151 => Ti := "010100011101111101100011001111011000000011001100"; --   +5365603   +4030668
      WHEN  152 => Ti := "010100100011111110011001001111001111111111100101"; --   +5390233   +3997669
      WHEN  153 => Ti := "010100101001111100000101001111000111111001101000"; --   +5414661   +3964520
      WHEN  154 => Ti := "010100101111110110100101001110111111110001010110"; --   +5438885   +3931222
      WHEN  155 => Ti := "010100110101101101111000001110110111100110110000"; --   +5462904   +3897776
      WHEN  156 => Ti := "010100111011100001111110001110101111011001110110"; --   +5486718   +3864182
      WHEN  157 => Ti := "010101000001010010110101001110100111001010101100"; --   +5510325   +3830444
      WHEN  158 => Ti := "010101000111000000011100001110011110111001010001"; --   +5533724   +3796561
      WHEN  159 => Ti := "010101001100101010110011001110010110100101100111"; --   +5556915   +3762535
      WHEN  160 => Ti := "010101010010010001111001001110001110001111110000"; --   +5579897   +3728368
      WHEN  161 => Ti := "010101010111110101101101001110000101110111101100"; --   +5602669   +3694060
      WHEN  162 => Ti := "010101011101010110001110001101111101011101011101"; --   +5625230   +3659613
      WHEN  163 => Ti := "010101100010110011011011001101110101000001000100"; --   +5647579   +3625028
      WHEN  164 => Ti := "010101101000001101010011001101101100100010100011"; --   +5669715   +3590307
      WHEN  165 => Ti := "010101101101100011110110001101100100000001111011"; --   +5691638   +3555451
      WHEN  166 => Ti := "010101110010110111000011001101011011011111001101"; --   +5713347   +3520461
      WHEN  167 => Ti := "010101111000000110111000001101010010111010011010"; --   +5734840   +3485338
      WHEN  168 => Ti := "010101111101010011010110001101001010010011100100"; --   +5756118   +3450084
      WHEN  169 => Ti := "010110000010011100011011001101000001101010101100"; --   +5777179   +3414700
      WHEN  170 => Ti := "010110000111100010000110001100111000111111110100"; --   +5798022   +3379188
      WHEN  171 => Ti := "010110001100100100011000001100110000010010111100"; --   +5818648   +3343548
      WHEN  172 => Ti := "010110010001100011001110001100100111100100000111"; --   +5839054   +3307783
      WHEN  173 => Ti := "010110010110011110101000001100011110110011010101"; --   +5859240   +3271893
      WHEN  174 => Ti := "010110011011010110100110001100010110000000101000"; --   +5879206   +3235880
      WHEN  175 => Ti := "010110100000001011000110001100001101001100000001"; --   +5898950   +3199745
      WHEN  176 => Ti := "010110100100111100001000001100000100010101100001"; --   +5918472   +3163489
      WHEN  177 => Ti := "010110101001101001101100001011111011011101001010"; --   +5937772   +3127114
      WHEN  178 => Ti := "010110101110010011101111001011110010100010111110"; --   +5956847   +3090622
      WHEN  179 => Ti := "010110110010111010010011001011101001100110111101"; --   +5975699   +3054013
      WHEN  180 => Ti := "010110110111011101010110001011100000101001001010"; --   +5994326   +3017290
      WHEN  181 => Ti := "010110111011111100110111001011010111101001100100"; --   +6012727   +2980452
      WHEN  182 => Ti := "010111000000011000110101001011001110101000001111"; --   +6030901   +2943503
      WHEN  183 => Ti := "010111000100110001010000001011000101100101001011"; --   +6048848   +2906443
      WHEN  184 => Ti := "010111001001000110001000001010111100100000011001"; --   +6066568   +2869273
      WHEN  185 => Ti := "010111001101010111011100001010110011011001111011"; --   +6084060   +2831995
      WHEN  186 => Ti := "010111010001100101001010001010101010010001110011"; --   +6101322   +2794611
      WHEN  187 => Ti := "010111010101101111010010001010100001001000000001"; --   +6118354   +2757121
      WHEN  188 => Ti := "010111011001110101110101001010010111111100101000"; --   +6135157   +2719528
      WHEN  189 => Ti := "010111011101111000110000001010001110101111101000"; --   +6151728   +2681832
      WHEN  190 => Ti := "010111100001111000000011001010000101100001000011"; --   +6168067   +2644035
      WHEN  191 => Ti := "010111100101110011101111001001111100010000111011"; --   +6184175   +2606139
      WHEN  192 => Ti := "010111101001101011110001001001110010111111010000"; --   +6200049   +2568144
      WHEN  193 => Ti := "010111101101100000001010001001101001101100000101"; --   +6215690   +2530053
      WHEN  194 => Ti := "010111110001010000111010001001100000010111011011"; --   +6231098   +2491867
      WHEN  195 => Ti := "010111110100111101111110001001010111000001010011"; --   +6246270   +2453587
      WHEN  196 => Ti := "010111111000100111010111001001001101101001101110"; --   +6261207   +2415214
      WHEN  197 => Ti := "010111111100001101000101001001000100010000101110"; --   +6275909   +2376750
      WHEN  198 => Ti := "010111111111101111000110001000111010110110010101"; --   +6290374   +2338197
      WHEN  199 => Ti := "011000000011001101011011001000110001011010100100"; --   +6304603   +2299556
      WHEN  200 => Ti := "011000000110101000000010001000100111111101011101"; --   +6318594   +2260829
      WHEN  201 => Ti := "011000001001111110111011001000011110011111000000"; --   +6332347   +2222016
      WHEN  202 => Ti := "011000001101010010000110001000010100111111010000"; --   +6345862   +2183120
      WHEN  203 => Ti := "011000010000100001100010001000001011011110001101"; --   +6359138   +2144141
      WHEN  204 => Ti := "011000010011101101001110001000000001111011111010"; --   +6372174   +2105082
      WHEN  205 => Ti := "011000010110110101001011000111111000011000010111"; --   +6384971   +2065943
      WHEN  206 => Ti := "011000011001111001010111000111101110110011100111"; --   +6397527   +2026727
      WHEN  207 => Ti := "011000011100111001110011000111100101001101101010"; --   +6409843   +1987434
      WHEN  208 => Ti := "011000011111110110011101000111011011100110100011"; --   +6421917   +1948067
      WHEN  209 => Ti := "011000100010101111010101000111010001111110010010"; --   +6433749   +1908626
      WHEN  210 => Ti := "011000100101100100011011000111001000010100111001"; --   +6445339   +1869113
      WHEN  211 => Ti := "011000101000010101101110000110111110101010011010"; --   +6456686   +1829530
      WHEN  212 => Ti := "011000101011000011001110000110110100111110110110"; --   +6467790   +1789878
      WHEN  213 => Ti := "011000101101101100111011000110101011010010001111"; --   +6478651   +1750159
      WHEN  214 => Ti := "011000110000010010110100000110100001100100100110"; --   +6489268   +1710374
      WHEN  215 => Ti := "011000110010110100111000000110010111110101111100"; --   +6499640   +1670524
      WHEN  216 => Ti := "011000110101010011001000000110001110000110010100"; --   +6509768   +1630612
      WHEN  217 => Ti := "011000110111101101100011000110000100010101101110"; --   +6519651   +1590638
      WHEN  218 => Ti := "011000111010000100001000000101111010100100001100"; --   +6529288   +1550604
      WHEN  219 => Ti := "011000111100010110111000000101110000110001110000"; --   +6538680   +1510512
      WHEN  220 => Ti := "011000111110100101110001000101100110111110011011"; --   +6547825   +1470363
      WHEN  221 => Ti := "011001000000110000110100000101011101001010001110"; --   +6556724   +1430158
      WHEN  222 => Ti := "011001000010110111111111000101010011010101001100"; --   +6565375   +1389900
      WHEN  223 => Ti := "011001000100111011010100000101001001011111010110"; --   +6573780   +1349590
      WHEN  224 => Ti := "011001000110111010110001000100111111101000101100"; --   +6581937   +1309228
      WHEN  225 => Ti := "011001001000110110010111000100110101110001010010"; --   +6589847   +1268818
      WHEN  226 => Ti := "011001001010101110000100000100101011111001000111"; --   +6597508   +1228359
      WHEN  227 => Ti := "011001001100100001111001000100100010000000001111"; --   +6604921   +1187855
      WHEN  228 => Ti := "011001001110010001110101000100011000000110101001"; --   +6612085   +1147305
      WHEN  229 => Ti := "011001001111111101111000000100001110001100011001"; --   +6619000   +1106713
      WHEN  230 => Ti := "011001010001100110000010000100000100010001011110"; --   +6625666   +1066078
      WHEN  231 => Ti := "011001010011001010010011000011111010010101111100"; --   +6632083   +1025404
      WHEN  232 => Ti := "011001010100101010101010000011110000011001110011"; --   +6638250    +984691
      WHEN  233 => Ti := "011001010110000111000111000011100110011101000101"; --   +6644167    +943941
      WHEN  234 => Ti := "011001010111011111101010000011011100011111110011"; --   +6649834    +903155
      WHEN  235 => Ti := "011001011000110100010010000011010010100010000000"; --   +6655250    +862336
      WHEN  236 => Ti := "011001011010000101000000000011001000100011101100"; --   +6660416    +821484
      WHEN  237 => Ti := "011001011011010001110011000010111110100100111001"; --   +6665331    +780601
      WHEN  238 => Ti := "011001011100011010101011000010110100100101101000"; --   +6669995    +739688
      WHEN  239 => Ti := "011001011101011111101001000010101010100101111100"; --   +6674409    +698748
      WHEN  240 => Ti := "011001011110100000101010000010100000100101110101"; --   +6678570    +657781
      WHEN  241 => Ti := "011001011111011101110001000010010110100101010110"; --   +6682481    +616790
      WHEN  242 => Ti := "011001100000010110111011000010001100100100011111"; --   +6686139    +575775
      WHEN  243 => Ti := "011001100001001100001010000010000010100011010011"; --   +6689546    +534739
      WHEN  244 => Ti := "011001100001111101011110000001111000100001110011"; --   +6692702    +493683
      WHEN  245 => Ti := "011001100010101010110101000001101110100000000000"; --   +6695605    +452608
      WHEN  246 => Ti := "011001100011010100010000000001100100011101111100"; --   +6698256    +411516
      WHEN  247 => Ti := "011001100011111001101111000001011010011011101000"; --   +6700655    +370408
      WHEN  248 => Ti := "011001100100011011010010000001010000011001000111"; --   +6702802    +329287
      WHEN  249 => Ti := "011001100100111000111000000001000110010110011001"; --   +6704696    +288153
      WHEN  250 => Ti := "011001100101010010100010000000111100010011100001"; --   +6706338    +247009
      WHEN  251 => Ti := "011001100101101000001111000000110010010000011111"; --   +6707727    +205855
      WHEN  252 => Ti := "011001100101111010000000000000101000001101010101"; --   +6708864    +164693
      WHEN  253 => Ti := "011001100110000111110100000000011110001010000101"; --   +6709748    +123525
      WHEN  254 => Ti := "011001100110010001101100000000010100000110110000"; --   +6710380     +82352
      WHEN  255 => Ti := "011001100110010111100111000000001010000011011001"; --   +6710759     +41177
      WHEN  256 => Ti := "011001100110011001100101000000000000000000000000"; --   +6710885         +0
      WHEN  257 => Ti := "011001100110010111100111111111110101111100100111"; --   +6710759     -41177
      WHEN  258 => Ti := "011001100110010001101100111111101011111001010000"; --   +6710380     -82352
      WHEN  259 => Ti := "011001100110000111110100111111100001110101111011"; --   +6709748    -123525
      WHEN  260 => Ti := "011001100101111010000000111111010111110010101011"; --   +6708864    -164693
      WHEN  261 => Ti := "011001100101101000001111111111001101101111100001"; --   +6707727    -205855
      WHEN  262 => Ti := "011001100101010010100010111111000011101100011111"; --   +6706338    -247009
      WHEN  263 => Ti := "011001100100111000111000111110111001101001100111"; --   +6704696    -288153
      WHEN  264 => Ti := "011001100100011011010010111110101111100110111001"; --   +6702802    -329287
      WHEN  265 => Ti := "011001100011111001101111111110100101100100011000"; --   +6700655    -370408
      WHEN  266 => Ti := "011001100011010100010000111110011011100010000100"; --   +6698256    -411516
      WHEN  267 => Ti := "011001100010101010110101111110010001100000000000"; --   +6695605    -452608
      WHEN  268 => Ti := "011001100001111101011110111110000111011110001101"; --   +6692702    -493683
      WHEN  269 => Ti := "011001100001001100001010111101111101011100101101"; --   +6689546    -534739
      WHEN  270 => Ti := "011001100000010110111011111101110011011011100001"; --   +6686139    -575775
      WHEN  271 => Ti := "011001011111011101110001111101101001011010101010"; --   +6682481    -616790
      WHEN  272 => Ti := "011001011110100000101010111101011111011010001011"; --   +6678570    -657781
      WHEN  273 => Ti := "011001011101011111101001111101010101011010000100"; --   +6674409    -698748
      WHEN  274 => Ti := "011001011100011010101011111101001011011010011000"; --   +6669995    -739688
      WHEN  275 => Ti := "011001011011010001110011111101000001011011000111"; --   +6665331    -780601
      WHEN  276 => Ti := "011001011010000101000000111100110111011100010100"; --   +6660416    -821484
      WHEN  277 => Ti := "011001011000110100010010111100101101011110000000"; --   +6655250    -862336
      WHEN  278 => Ti := "011001010111011111101010111100100011100000001101"; --   +6649834    -903155
      WHEN  279 => Ti := "011001010110000111000111111100011001100010111011"; --   +6644167    -943941
      WHEN  280 => Ti := "011001010100101010101010111100001111100110001101"; --   +6638250    -984691
      WHEN  281 => Ti := "011001010011001010010011111100000101101010000100"; --   +6632083   -1025404
      WHEN  282 => Ti := "011001010001100110000010111011111011101110100010"; --   +6625666   -1066078
      WHEN  283 => Ti := "011001001111111101111000111011110001110011100111"; --   +6619000   -1106713
      WHEN  284 => Ti := "011001001110010001110101111011100111111001010111"; --   +6612085   -1147305
      WHEN  285 => Ti := "011001001100100001111001111011011101111111110001"; --   +6604921   -1187855
      WHEN  286 => Ti := "011001001010101110000100111011010100000110111001"; --   +6597508   -1228359
      WHEN  287 => Ti := "011001001000110110010111111011001010001110101110"; --   +6589847   -1268818
      WHEN  288 => Ti := "011001000110111010110001111011000000010111010100"; --   +6581937   -1309228
      WHEN  289 => Ti := "011001000100111011010100111010110110100000101010"; --   +6573780   -1349590
      WHEN  290 => Ti := "011001000010110111111111111010101100101010110100"; --   +6565375   -1389900
      WHEN  291 => Ti := "011001000000110000110100111010100010110101110010"; --   +6556724   -1430158
      WHEN  292 => Ti := "011000111110100101110001111010011001000001100101"; --   +6547825   -1470363
      WHEN  293 => Ti := "011000111100010110111000111010001111001110010000"; --   +6538680   -1510512
      WHEN  294 => Ti := "011000111010000100001000111010000101011011110100"; --   +6529288   -1550604
      WHEN  295 => Ti := "011000110111101101100011111001111011101010010010"; --   +6519651   -1590638
      WHEN  296 => Ti := "011000110101010011001000111001110001111001101100"; --   +6509768   -1630612
      WHEN  297 => Ti := "011000110010110100111000111001101000001010000100"; --   +6499640   -1670524
      WHEN  298 => Ti := "011000110000010010110100111001011110011011011010"; --   +6489268   -1710374
      WHEN  299 => Ti := "011000101101101100111011111001010100101101110001"; --   +6478651   -1750159
      WHEN  300 => Ti := "011000101011000011001110111001001011000001001010"; --   +6467790   -1789878
      WHEN  301 => Ti := "011000101000010101101110111001000001010101100110"; --   +6456686   -1829530
      WHEN  302 => Ti := "011000100101100100011011111000110111101011000111"; --   +6445339   -1869113
      WHEN  303 => Ti := "011000100010101111010101111000101110000001101110"; --   +6433749   -1908626
      WHEN  304 => Ti := "011000011111110110011101111000100100011001011101"; --   +6421917   -1948067
      WHEN  305 => Ti := "011000011100111001110011111000011010110010010110"; --   +6409843   -1987434
      WHEN  306 => Ti := "011000011001111001010111111000010001001100011001"; --   +6397527   -2026727
      WHEN  307 => Ti := "011000010110110101001011111000000111100111101001"; --   +6384971   -2065943
      WHEN  308 => Ti := "011000010011101101001110110111111110000100000110"; --   +6372174   -2105082
      WHEN  309 => Ti := "011000010000100001100010110111110100100001110011"; --   +6359138   -2144141
      WHEN  310 => Ti := "011000001101010010000110110111101011000000110000"; --   +6345862   -2183120
      WHEN  311 => Ti := "011000001001111110111011110111100001100001000000"; --   +6332347   -2222016
      WHEN  312 => Ti := "011000000110101000000010110111011000000010100011"; --   +6318594   -2260829
      WHEN  313 => Ti := "011000000011001101011011110111001110100101011100"; --   +6304603   -2299556
      WHEN  314 => Ti := "010111111111101111000110110111000101001001101011"; --   +6290374   -2338197
      WHEN  315 => Ti := "010111111100001101000101110110111011101111010010"; --   +6275909   -2376750
      WHEN  316 => Ti := "010111111000100111010111110110110010010110010010"; --   +6261207   -2415214
      WHEN  317 => Ti := "010111110100111101111110110110101000111110101101"; --   +6246270   -2453587
      WHEN  318 => Ti := "010111110001010000111010110110011111101000100101"; --   +6231098   -2491867
      WHEN  319 => Ti := "010111101101100000001010110110010110010011111011"; --   +6215690   -2530053
      WHEN  320 => Ti := "010111101001101011110001110110001101000000110000"; --   +6200049   -2568144
      WHEN  321 => Ti := "010111100101110011101111110110000011101111000101"; --   +6184175   -2606139
      WHEN  322 => Ti := "010111100001111000000011110101111010011110111101"; --   +6168067   -2644035
      WHEN  323 => Ti := "010111011101111000110000110101110001010000011000"; --   +6151728   -2681832
      WHEN  324 => Ti := "010111011001110101110101110101101000000011011000"; --   +6135157   -2719528
      WHEN  325 => Ti := "010111010101101111010010110101011110110111111111"; --   +6118354   -2757121
      WHEN  326 => Ti := "010111010001100101001010110101010101101110001101"; --   +6101322   -2794611
      WHEN  327 => Ti := "010111001101010111011100110101001100100110000101"; --   +6084060   -2831995
      WHEN  328 => Ti := "010111001001000110001000110101000011011111100111"; --   +6066568   -2869273
      WHEN  329 => Ti := "010111000100110001010000110100111010011010110101"; --   +6048848   -2906443
      WHEN  330 => Ti := "010111000000011000110101110100110001010111110001"; --   +6030901   -2943503
      WHEN  331 => Ti := "010110111011111100110111110100101000010110011100"; --   +6012727   -2980452
      WHEN  332 => Ti := "010110110111011101010110110100011111010110110110"; --   +5994326   -3017290
      WHEN  333 => Ti := "010110110010111010010011110100010110011001000011"; --   +5975699   -3054013
      WHEN  334 => Ti := "010110101110010011101111110100001101011101000010"; --   +5956847   -3090622
      WHEN  335 => Ti := "010110101001101001101100110100000100100010110110"; --   +5937772   -3127114
      WHEN  336 => Ti := "010110100100111100001000110011111011101010011111"; --   +5918472   -3163489
      WHEN  337 => Ti := "010110100000001011000110110011110010110011111111"; --   +5898950   -3199745
      WHEN  338 => Ti := "010110011011010110100110110011101001111111011000"; --   +5879206   -3235880
      WHEN  339 => Ti := "010110010110011110101000110011100001001100101011"; --   +5859240   -3271893
      WHEN  340 => Ti := "010110010001100011001110110011011000011011111001"; --   +5839054   -3307783
      WHEN  341 => Ti := "010110001100100100011000110011001111101101000100"; --   +5818648   -3343548
      WHEN  342 => Ti := "010110000111100010000110110011000111000000001100"; --   +5798022   -3379188
      WHEN  343 => Ti := "010110000010011100011011110010111110010101010100"; --   +5777179   -3414700
      WHEN  344 => Ti := "010101111101010011010110110010110101101100011100"; --   +5756118   -3450084
      WHEN  345 => Ti := "010101111000000110111000110010101101000101100110"; --   +5734840   -3485338
      WHEN  346 => Ti := "010101110010110111000011110010100100100000110011"; --   +5713347   -3520461
      WHEN  347 => Ti := "010101101101100011110110110010011011111110000101"; --   +5691638   -3555451
      WHEN  348 => Ti := "010101101000001101010011110010010011011101011101"; --   +5669715   -3590307
      WHEN  349 => Ti := "010101100010110011011011110010001010111110111100"; --   +5647579   -3625028
      WHEN  350 => Ti := "010101011101010110001110110010000010100010100011"; --   +5625230   -3659613
      WHEN  351 => Ti := "010101010111110101101101110001111010001000010100"; --   +5602669   -3694060
      WHEN  352 => Ti := "010101010010010001111001110001110001110000010000"; --   +5579897   -3728368
      WHEN  353 => Ti := "010101001100101010110011110001101001011010011001"; --   +5556915   -3762535
      WHEN  354 => Ti := "010101000111000000011100110001100001000110101111"; --   +5533724   -3796561
      WHEN  355 => Ti := "010101000001010010110101110001011000110101010100"; --   +5510325   -3830444
      WHEN  356 => Ti := "010100111011100001111110110001010000100110001010"; --   +5486718   -3864182
      WHEN  357 => Ti := "010100110101101101111000110001001000011001010000"; --   +5462904   -3897776
      WHEN  358 => Ti := "010100101111110110100101110001000000001110101010"; --   +5438885   -3931222
      WHEN  359 => Ti := "010100101001111100000101110000111000000110011000"; --   +5414661   -3964520
      WHEN  360 => Ti := "010100100011111110011001110000110000000000011011"; --   +5390233   -3997669
      WHEN  361 => Ti := "010100011101111101100011110000100111111100110100"; --   +5365603   -4030668
      WHEN  362 => Ti := "010100010111111001100010110000011111111011100101"; --   +5340770   -4063515
      WHEN  363 => Ti := "010100010001110010011000110000010111111100101111"; --   +5315736   -4096209
      WHEN  364 => Ti := "010100001011101000000110110000010000000000010100"; --   +5290502   -4128748
      WHEN  365 => Ti := "010100000101011010101101110000001000000110010011"; --   +5265069   -4161133
      WHEN  366 => Ti := "010011111111001010001110110000000000001110110000"; --   +5239438   -4193360
      WHEN  367 => Ti := "010011111000110110101001101111111000011001101010"; --   +5213609   -4225430
      WHEN  368 => Ti := "010011110010100000000000101111110000100111000100"; --   +5187584   -4257340
      WHEN  369 => Ti := "010011101100000110010100101111101000110110111101"; --   +5161364   -4289091
      WHEN  370 => Ti := "010011100101101001100101101111100001001001011001"; --   +5134949   -4320679
      WHEN  371 => Ti := "010011011111001001110110101111011001011110010111"; --   +5108342   -4352105
      WHEN  372 => Ti := "010011011000100111000101101111010001110101111000"; --   +5081541   -4383368
      WHEN  373 => Ti := "010011010010000001010110101111001010001111111111"; --   +5054550   -4414465
      WHEN  374 => Ti := "010011001011011000101000101111000010101100101100"; --   +5027368   -4445396
      WHEN  375 => Ti := "010011000100101100111101101110111011001100000000"; --   +4999997   -4476160
      WHEN  376 => Ti := "010010111101111110010110101110110011101101111101"; --   +4972438   -4506755
      WHEN  377 => Ti := "010010110111001100110011101110101100010010100100"; --   +4944691   -4537180
      WHEN  378 => Ti := "010010110000011000010111101110100100111001110101"; --   +4916759   -4567435
      WHEN  379 => Ti := "010010101001100001000001101110011101100011110010"; --   +4888641   -4597518
      WHEN  380 => Ti := "010010100010100110110011101110010110010000011101"; --   +4860339   -4627427
      WHEN  381 => Ti := "010010011011101001101110101110001110111111110101"; --   +4831854   -4657163
      WHEN  382 => Ti := "010010010100101001110011101110000111110001111101"; --   +4803187   -4686723
      WHEN  383 => Ti := "010010001101100111000100101110000000100110110110"; --   +4774340   -4716106
      WHEN  384 => Ti := "010010000110100001100000101101111001011110100000"; --   +4745312   -4745312
      WHEN  385 => Ti := "010001111111011001001010101101110010011000111100"; --   +4716106   -4774340
      WHEN  386 => Ti := "010001111000001110000011101101101011010110001101"; --   +4686723   -4803187
      WHEN  387 => Ti := "010001110001000000001011101101100100010110010010"; --   +4657163   -4831854
      WHEN  388 => Ti := "010001101001101111100011101101011101011001001101"; --   +4627427   -4860339
      WHEN  389 => Ti := "010001100010011100001110101101010110011110111111"; --   +4597518   -4888641
      WHEN  390 => Ti := "010001011011000110001011101101001111100111101001"; --   +4567435   -4916759
      WHEN  391 => Ti := "010001010011101101011100101101001000110011001101"; --   +4537180   -4944691
      WHEN  392 => Ti := "010001001100010010000011101101000010000001101010"; --   +4506755   -4972438
      WHEN  393 => Ti := "010001000100110100000000101100111011010011000011"; --   +4476160   -4999997
      WHEN  394 => Ti := "010000111101010011010100101100110100100111011000"; --   +4445396   -5027368
      WHEN  395 => Ti := "010000110101110000000001101100101101111110101010"; --   +4414465   -5054550
      WHEN  396 => Ti := "010000101110001010001000101100100111011000111011"; --   +4383368   -5081541
      WHEN  397 => Ti := "010000100110100001101001101100100000110110001010"; --   +4352105   -5108342
      WHEN  398 => Ti := "010000011110110110100111101100011010010110011011"; --   +4320679   -5134949
      WHEN  399 => Ti := "010000010111001001000011101100010011111001101100"; --   +4289091   -5161364
      WHEN  400 => Ti := "010000001111011000111100101100001101100000000000"; --   +4257340   -5187584
      WHEN  401 => Ti := "010000000111100110010110101100000111001001010111"; --   +4225430   -5213609
      WHEN  402 => Ti := "001111111111110001010000101100000000110101110010"; --   +4193360   -5239438
      WHEN  403 => Ti := "001111110111111001101101101011111010100101010011"; --   +4161133   -5265069
      WHEN  404 => Ti := "001111101111111111101100101011110100010111111010"; --   +4128748   -5290502
      WHEN  405 => Ti := "001111101000000011010001101011101110001101101000"; --   +4096209   -5315736
      WHEN  406 => Ti := "001111100000000100011011101011101000000110011110"; --   +4063515   -5340770
      WHEN  407 => Ti := "001111011000000011001100101011100010000010011101"; --   +4030668   -5365603
      WHEN  408 => Ti := "001111001111111111100101101011011100000001100111"; --   +3997669   -5390233
      WHEN  409 => Ti := "001111000111111001101000101011010110000011111011"; --   +3964520   -5414661
      WHEN  410 => Ti := "001110111111110001010110101011010000001001011011"; --   +3931222   -5438885
      WHEN  411 => Ti := "001110110111100110110000101011001010010010001000"; --   +3897776   -5462904
      WHEN  412 => Ti := "001110101111011001110110101011000100011110000010"; --   +3864182   -5486718
      WHEN  413 => Ti := "001110100111001010101100101010111110101101001011"; --   +3830444   -5510325
      WHEN  414 => Ti := "001110011110111001010001101010111000111111100100"; --   +3796561   -5533724
      WHEN  415 => Ti := "001110010110100101100111101010110011010101001101"; --   +3762535   -5556915
      WHEN  416 => Ti := "001110001110001111110000101010101101101110000111"; --   +3728368   -5579897
      WHEN  417 => Ti := "001110000101110111101100101010101000001010010011"; --   +3694060   -5602669
      WHEN  418 => Ti := "001101111101011101011101101010100010101001110010"; --   +3659613   -5625230
      WHEN  419 => Ti := "001101110101000001000100101010011101001100100101"; --   +3625028   -5647579
      WHEN  420 => Ti := "001101101100100010100011101010010111110010101101"; --   +3590307   -5669715
      WHEN  421 => Ti := "001101100100000001111011101010010010011100001010"; --   +3555451   -5691638
      WHEN  422 => Ti := "001101011011011111001101101010001101001000111101"; --   +3520461   -5713347
      WHEN  423 => Ti := "001101010010111010011010101010000111111001001000"; --   +3485338   -5734840
      WHEN  424 => Ti := "001101001010010011100100101010000010101100101010"; --   +3450084   -5756118
      WHEN  425 => Ti := "001101000001101010101100101001111101100011100101"; --   +3414700   -5777179
      WHEN  426 => Ti := "001100111000111111110100101001111000011101111010"; --   +3379188   -5798022
      WHEN  427 => Ti := "001100110000010010111100101001110011011011101000"; --   +3343548   -5818648
      WHEN  428 => Ti := "001100100111100100000111101001101110011100110010"; --   +3307783   -5839054
      WHEN  429 => Ti := "001100011110110011010101101001101001100001011000"; --   +3271893   -5859240
      WHEN  430 => Ti := "001100010110000000101000101001100100101001011010"; --   +3235880   -5879206
      WHEN  431 => Ti := "001100001101001100000001101001011111110100111010"; --   +3199745   -5898950
      WHEN  432 => Ti := "001100000100010101100001101001011011000011111000"; --   +3163489   -5918472
      WHEN  433 => Ti := "001011111011011101001010101001010110010110010100"; --   +3127114   -5937772
      WHEN  434 => Ti := "001011110010100010111110101001010001101100010001"; --   +3090622   -5956847
      WHEN  435 => Ti := "001011101001100110111101101001001101000101101101"; --   +3054013   -5975699
      WHEN  436 => Ti := "001011100000101001001010101001001000100010101010"; --   +3017290   -5994326
      WHEN  437 => Ti := "001011010111101001100100101001000100000011001001"; --   +2980452   -6012727
      WHEN  438 => Ti := "001011001110101000001111101000111111100111001011"; --   +2943503   -6030901
      WHEN  439 => Ti := "001011000101100101001011101000111011001110110000"; --   +2906443   -6048848
      WHEN  440 => Ti := "001010111100100000011001101000110110111001111000"; --   +2869273   -6066568
      WHEN  441 => Ti := "001010110011011001111011101000110010101000100100"; --   +2831995   -6084060
      WHEN  442 => Ti := "001010101010010001110011101000101110011010110110"; --   +2794611   -6101322
      WHEN  443 => Ti := "001010100001001000000001101000101010010000101110"; --   +2757121   -6118354
      WHEN  444 => Ti := "001010010111111100101000101000100110001010001011"; --   +2719528   -6135157
      WHEN  445 => Ti := "001010001110101111101000101000100010000111010000"; --   +2681832   -6151728
      WHEN  446 => Ti := "001010000101100001000011101000011110000111111101"; --   +2644035   -6168067
      WHEN  447 => Ti := "001001111100010000111011101000011010001100010001"; --   +2606139   -6184175
      WHEN  448 => Ti := "001001110010111111010000101000010110010100001111"; --   +2568144   -6200049
      WHEN  449 => Ti := "001001101001101100000101101000010010011111110110"; --   +2530053   -6215690
      WHEN  450 => Ti := "001001100000010111011011101000001110101111000110"; --   +2491867   -6231098
      WHEN  451 => Ti := "001001010111000001010011101000001011000010000010"; --   +2453587   -6246270
      WHEN  452 => Ti := "001001001101101001101110101000000111011000101001"; --   +2415214   -6261207
      WHEN  453 => Ti := "001001000100010000101110101000000011110010111011"; --   +2376750   -6275909
      WHEN  454 => Ti := "001000111010110110010101101000000000010000111010"; --   +2338197   -6290374
      WHEN  455 => Ti := "001000110001011010100100100111111100110010100101"; --   +2299556   -6304603
      WHEN  456 => Ti := "001000100111111101011101100111111001010111111110"; --   +2260829   -6318594
      WHEN  457 => Ti := "001000011110011111000000100111110110000001000101"; --   +2222016   -6332347
      WHEN  458 => Ti := "001000010100111111010000100111110010101101111010"; --   +2183120   -6345862
      WHEN  459 => Ti := "001000001011011110001101100111101111011110011110"; --   +2144141   -6359138
      WHEN  460 => Ti := "001000000001111011111010100111101100010010110010"; --   +2105082   -6372174
      WHEN  461 => Ti := "000111111000011000010111100111101001001010110101"; --   +2065943   -6384971
      WHEN  462 => Ti := "000111101110110011100111100111100110000110101001"; --   +2026727   -6397527
      WHEN  463 => Ti := "000111100101001101101010100111100011000110001101"; --   +1987434   -6409843
      WHEN  464 => Ti := "000111011011100110100011100111100000001001100011"; --   +1948067   -6421917
      WHEN  465 => Ti := "000111010001111110010010100111011101010000101011"; --   +1908626   -6433749
      WHEN  466 => Ti := "000111001000010100111001100111011010011011100101"; --   +1869113   -6445339
      WHEN  467 => Ti := "000110111110101010011010100111010111101010010010"; --   +1829530   -6456686
      WHEN  468 => Ti := "000110110100111110110110100111010100111100110010"; --   +1789878   -6467790
      WHEN  469 => Ti := "000110101011010010001111100111010010010011000101"; --   +1750159   -6478651
      WHEN  470 => Ti := "000110100001100100100110100111001111101101001100"; --   +1710374   -6489268
      WHEN  471 => Ti := "000110010111110101111100100111001101001011001000"; --   +1670524   -6499640
      WHEN  472 => Ti := "000110001110000110010100100111001010101100111000"; --   +1630612   -6509768
      WHEN  473 => Ti := "000110000100010101101110100111001000010010011101"; --   +1590638   -6519651
      WHEN  474 => Ti := "000101111010100100001100100111000101111011111000"; --   +1550604   -6529288
      WHEN  475 => Ti := "000101110000110001110000100111000011101001001000"; --   +1510512   -6538680
      WHEN  476 => Ti := "000101100110111110011011100111000001011010001111"; --   +1470363   -6547825
      WHEN  477 => Ti := "000101011101001010001110100110111111001111001100"; --   +1430158   -6556724
      WHEN  478 => Ti := "000101010011010101001100100110111101001000000001"; --   +1389900   -6565375
      WHEN  479 => Ti := "000101001001011111010110100110111011000100101100"; --   +1349590   -6573780
      WHEN  480 => Ti := "000100111111101000101100100110111001000101001111"; --   +1309228   -6581937
      WHEN  481 => Ti := "000100110101110001010010100110110111001001101001"; --   +1268818   -6589847
      WHEN  482 => Ti := "000100101011111001000111100110110101010001111100"; --   +1228359   -6597508
      WHEN  483 => Ti := "000100100010000000001111100110110011011110000111"; --   +1187855   -6604921
      WHEN  484 => Ti := "000100011000000110101001100110110001101110001011"; --   +1147305   -6612085
      WHEN  485 => Ti := "000100001110001100011001100110110000000010001000"; --   +1106713   -6619000
      WHEN  486 => Ti := "000100000100010001011110100110101110011001111110"; --   +1066078   -6625666
      WHEN  487 => Ti := "000011111010010101111100100110101100110101101101"; --   +1025404   -6632083
      WHEN  488 => Ti := "000011110000011001110011100110101011010101010110"; --    +984691   -6638250
      WHEN  489 => Ti := "000011100110011101000101100110101001111000111001"; --    +943941   -6644167
      WHEN  490 => Ti := "000011011100011111110011100110101000100000010110"; --    +903155   -6649834
      WHEN  491 => Ti := "000011010010100010000000100110100111001011101110"; --    +862336   -6655250
      WHEN  492 => Ti := "000011001000100011101100100110100101111011000000"; --    +821484   -6660416
      WHEN  493 => Ti := "000010111110100100111001100110100100101110001101"; --    +780601   -6665331
      WHEN  494 => Ti := "000010110100100101101000100110100011100101010101"; --    +739688   -6669995
      WHEN  495 => Ti := "000010101010100101111100100110100010100000010111"; --    +698748   -6674409
      WHEN  496 => Ti := "000010100000100101110101100110100001011111010110"; --    +657781   -6678570
      WHEN  497 => Ti := "000010010110100101010110100110100000100010001111"; --    +616790   -6682481
      WHEN  498 => Ti := "000010001100100100011111100110011111101001000101"; --    +575775   -6686139
      WHEN  499 => Ti := "000010000010100011010011100110011110110011110110"; --    +534739   -6689546
      WHEN  500 => Ti := "000001111000100001110011100110011110000010100010"; --    +493683   -6692702
      WHEN  501 => Ti := "000001101110100000000000100110011101010101001011"; --    +452608   -6695605
      WHEN  502 => Ti := "000001100100011101111100100110011100101011110000"; --    +411516   -6698256
      WHEN  503 => Ti := "000001011010011011101000100110011100000110010001"; --    +370408   -6700655
      WHEN  504 => Ti := "000001010000011001000111100110011011100100101110"; --    +329287   -6702802
      WHEN  505 => Ti := "000001000110010110011001100110011011000111001000"; --    +288153   -6704696
      WHEN  506 => Ti := "000000111100010011100001100110011010101101011110"; --    +247009   -6706338
      WHEN  507 => Ti := "000000110010010000011111100110011010010111110001"; --    +205855   -6707727
      WHEN  508 => Ti := "000000101000001101010101100110011010000110000000"; --    +164693   -6708864
      WHEN  509 => Ti := "000000011110001010000101100110011001111000001100"; --    +123525   -6709748
      WHEN  510 => Ti := "000000010100000110110000100110011001101110010100"; --     +82352   -6710380
      WHEN  511 => Ti := "000000001010000011011001100110011001101000011001"; --     +41177   -6710759
      WHEN  512 => Ti := "000000000000000000000000100110011001100110011011"; --         +0   -6710885
      WHEN  513 => Ti := "111111110101111100100111100110011001101000011001"; --     -41177   -6710759
      WHEN  514 => Ti := "111111101011111001010000100110011001101110010100"; --     -82352   -6710380
      WHEN  515 => Ti := "111111100001110101111011100110011001111000001100"; --    -123525   -6709748
      WHEN  516 => Ti := "111111010111110010101011100110011010000110000000"; --    -164693   -6708864
      WHEN  517 => Ti := "111111001101101111100001100110011010010111110001"; --    -205855   -6707727
      WHEN  518 => Ti := "111111000011101100011111100110011010101101011110"; --    -247009   -6706338
      WHEN  519 => Ti := "111110111001101001100111100110011011000111001000"; --    -288153   -6704696
      WHEN  520 => Ti := "111110101111100110111001100110011011100100101110"; --    -329287   -6702802
      WHEN  521 => Ti := "111110100101100100011000100110011100000110010001"; --    -370408   -6700655
      WHEN  522 => Ti := "111110011011100010000100100110011100101011110000"; --    -411516   -6698256
      WHEN  523 => Ti := "111110010001100000000000100110011101010101001011"; --    -452608   -6695605
      WHEN  524 => Ti := "111110000111011110001101100110011110000010100010"; --    -493683   -6692702
      WHEN  525 => Ti := "111101111101011100101101100110011110110011110110"; --    -534739   -6689546
      WHEN  526 => Ti := "111101110011011011100001100110011111101001000101"; --    -575775   -6686139
      WHEN  527 => Ti := "111101101001011010101010100110100000100010001111"; --    -616790   -6682481
      WHEN  528 => Ti := "111101011111011010001011100110100001011111010110"; --    -657781   -6678570
      WHEN  529 => Ti := "111101010101011010000100100110100010100000010111"; --    -698748   -6674409
      WHEN  530 => Ti := "111101001011011010011000100110100011100101010101"; --    -739688   -6669995
      WHEN  531 => Ti := "111101000001011011000111100110100100101110001101"; --    -780601   -6665331
      WHEN  532 => Ti := "111100110111011100010100100110100101111011000000"; --    -821484   -6660416
      WHEN  533 => Ti := "111100101101011110000000100110100111001011101110"; --    -862336   -6655250
      WHEN  534 => Ti := "111100100011100000001101100110101000100000010110"; --    -903155   -6649834
      WHEN  535 => Ti := "111100011001100010111011100110101001111000111001"; --    -943941   -6644167
      WHEN  536 => Ti := "111100001111100110001101100110101011010101010110"; --    -984691   -6638250
      WHEN  537 => Ti := "111100000101101010000100100110101100110101101101"; --   -1025404   -6632083
      WHEN  538 => Ti := "111011111011101110100010100110101110011001111110"; --   -1066078   -6625666
      WHEN  539 => Ti := "111011110001110011100111100110110000000010001000"; --   -1106713   -6619000
      WHEN  540 => Ti := "111011100111111001010111100110110001101110001011"; --   -1147305   -6612085
      WHEN  541 => Ti := "111011011101111111110001100110110011011110000111"; --   -1187855   -6604921
      WHEN  542 => Ti := "111011010100000110111001100110110101010001111100"; --   -1228359   -6597508
      WHEN  543 => Ti := "111011001010001110101110100110110111001001101001"; --   -1268818   -6589847
      WHEN  544 => Ti := "111011000000010111010100100110111001000101001111"; --   -1309228   -6581937
      WHEN  545 => Ti := "111010110110100000101010100110111011000100101100"; --   -1349590   -6573780
      WHEN  546 => Ti := "111010101100101010110100100110111101001000000001"; --   -1389900   -6565375
      WHEN  547 => Ti := "111010100010110101110010100110111111001111001100"; --   -1430158   -6556724
      WHEN  548 => Ti := "111010011001000001100101100111000001011010001111"; --   -1470363   -6547825
      WHEN  549 => Ti := "111010001111001110010000100111000011101001001000"; --   -1510512   -6538680
      WHEN  550 => Ti := "111010000101011011110100100111000101111011111000"; --   -1550604   -6529288
      WHEN  551 => Ti := "111001111011101010010010100111001000010010011101"; --   -1590638   -6519651
      WHEN  552 => Ti := "111001110001111001101100100111001010101100111000"; --   -1630612   -6509768
      WHEN  553 => Ti := "111001101000001010000100100111001101001011001000"; --   -1670524   -6499640
      WHEN  554 => Ti := "111001011110011011011010100111001111101101001100"; --   -1710374   -6489268
      WHEN  555 => Ti := "111001010100101101110001100111010010010011000101"; --   -1750159   -6478651
      WHEN  556 => Ti := "111001001011000001001010100111010100111100110010"; --   -1789878   -6467790
      WHEN  557 => Ti := "111001000001010101100110100111010111101010010010"; --   -1829530   -6456686
      WHEN  558 => Ti := "111000110111101011000111100111011010011011100101"; --   -1869113   -6445339
      WHEN  559 => Ti := "111000101110000001101110100111011101010000101011"; --   -1908626   -6433749
      WHEN  560 => Ti := "111000100100011001011101100111100000001001100011"; --   -1948067   -6421917
      WHEN  561 => Ti := "111000011010110010010110100111100011000110001101"; --   -1987434   -6409843
      WHEN  562 => Ti := "111000010001001100011001100111100110000110101001"; --   -2026727   -6397527
      WHEN  563 => Ti := "111000000111100111101001100111101001001010110101"; --   -2065943   -6384971
      WHEN  564 => Ti := "110111111110000100000110100111101100010010110010"; --   -2105082   -6372174
      WHEN  565 => Ti := "110111110100100001110011100111101111011110011110"; --   -2144141   -6359138
      WHEN  566 => Ti := "110111101011000000110000100111110010101101111010"; --   -2183120   -6345862
      WHEN  567 => Ti := "110111100001100001000000100111110110000001000101"; --   -2222016   -6332347
      WHEN  568 => Ti := "110111011000000010100011100111111001010111111110"; --   -2260829   -6318594
      WHEN  569 => Ti := "110111001110100101011100100111111100110010100101"; --   -2299556   -6304603
      WHEN  570 => Ti := "110111000101001001101011101000000000010000111010"; --   -2338197   -6290374
      WHEN  571 => Ti := "110110111011101111010010101000000011110010111011"; --   -2376750   -6275909
      WHEN  572 => Ti := "110110110010010110010010101000000111011000101001"; --   -2415214   -6261207
      WHEN  573 => Ti := "110110101000111110101101101000001011000010000010"; --   -2453587   -6246270
      WHEN  574 => Ti := "110110011111101000100101101000001110101111000110"; --   -2491867   -6231098
      WHEN  575 => Ti := "110110010110010011111011101000010010011111110110"; --   -2530053   -6215690
      WHEN  576 => Ti := "110110001101000000110000101000010110010100001111"; --   -2568144   -6200049
      WHEN  577 => Ti := "110110000011101111000101101000011010001100010001"; --   -2606139   -6184175
      WHEN  578 => Ti := "110101111010011110111101101000011110000111111101"; --   -2644035   -6168067
      WHEN  579 => Ti := "110101110001010000011000101000100010000111010000"; --   -2681832   -6151728
      WHEN  580 => Ti := "110101101000000011011000101000100110001010001011"; --   -2719528   -6135157
      WHEN  581 => Ti := "110101011110110111111111101000101010010000101110"; --   -2757121   -6118354
      WHEN  582 => Ti := "110101010101101110001101101000101110011010110110"; --   -2794611   -6101322
      WHEN  583 => Ti := "110101001100100110000101101000110010101000100100"; --   -2831995   -6084060
      WHEN  584 => Ti := "110101000011011111100111101000110110111001111000"; --   -2869273   -6066568
      WHEN  585 => Ti := "110100111010011010110101101000111011001110110000"; --   -2906443   -6048848
      WHEN  586 => Ti := "110100110001010111110001101000111111100111001011"; --   -2943503   -6030901
      WHEN  587 => Ti := "110100101000010110011100101001000100000011001001"; --   -2980452   -6012727
      WHEN  588 => Ti := "110100011111010110110110101001001000100010101010"; --   -3017290   -5994326
      WHEN  589 => Ti := "110100010110011001000011101001001101000101101101"; --   -3054013   -5975699
      WHEN  590 => Ti := "110100001101011101000010101001010001101100010001"; --   -3090622   -5956847
      WHEN  591 => Ti := "110100000100100010110110101001010110010110010100"; --   -3127114   -5937772
      WHEN  592 => Ti := "110011111011101010011111101001011011000011111000"; --   -3163489   -5918472
      WHEN  593 => Ti := "110011110010110011111111101001011111110100111010"; --   -3199745   -5898950
      WHEN  594 => Ti := "110011101001111111011000101001100100101001011010"; --   -3235880   -5879206
      WHEN  595 => Ti := "110011100001001100101011101001101001100001011000"; --   -3271893   -5859240
      WHEN  596 => Ti := "110011011000011011111001101001101110011100110010"; --   -3307783   -5839054
      WHEN  597 => Ti := "110011001111101101000100101001110011011011101000"; --   -3343548   -5818648
      WHEN  598 => Ti := "110011000111000000001100101001111000011101111010"; --   -3379188   -5798022
      WHEN  599 => Ti := "110010111110010101010100101001111101100011100101"; --   -3414700   -5777179
      WHEN  600 => Ti := "110010110101101100011100101010000010101100101010"; --   -3450084   -5756118
      WHEN  601 => Ti := "110010101101000101100110101010000111111001001000"; --   -3485338   -5734840
      WHEN  602 => Ti := "110010100100100000110011101010001101001000111101"; --   -3520461   -5713347
      WHEN  603 => Ti := "110010011011111110000101101010010010011100001010"; --   -3555451   -5691638
      WHEN  604 => Ti := "110010010011011101011101101010010111110010101101"; --   -3590307   -5669715
      WHEN  605 => Ti := "110010001010111110111100101010011101001100100101"; --   -3625028   -5647579
      WHEN  606 => Ti := "110010000010100010100011101010100010101001110010"; --   -3659613   -5625230
      WHEN  607 => Ti := "110001111010001000010100101010101000001010010011"; --   -3694060   -5602669
      WHEN  608 => Ti := "110001110001110000010000101010101101101110000111"; --   -3728368   -5579897
      WHEN  609 => Ti := "110001101001011010011001101010110011010101001101"; --   -3762535   -5556915
      WHEN  610 => Ti := "110001100001000110101111101010111000111111100100"; --   -3796561   -5533724
      WHEN  611 => Ti := "110001011000110101010100101010111110101101001011"; --   -3830444   -5510325
      WHEN  612 => Ti := "110001010000100110001010101011000100011110000010"; --   -3864182   -5486718
      WHEN  613 => Ti := "110001001000011001010000101011001010010010001000"; --   -3897776   -5462904
      WHEN  614 => Ti := "110001000000001110101010101011010000001001011011"; --   -3931222   -5438885
      WHEN  615 => Ti := "110000111000000110011000101011010110000011111011"; --   -3964520   -5414661
      WHEN  616 => Ti := "110000110000000000011011101011011100000001100111"; --   -3997669   -5390233
      WHEN  617 => Ti := "110000100111111100110100101011100010000010011101"; --   -4030668   -5365603
      WHEN  618 => Ti := "110000011111111011100101101011101000000110011110"; --   -4063515   -5340770
      WHEN  619 => Ti := "110000010111111100101111101011101110001101101000"; --   -4096209   -5315736
      WHEN  620 => Ti := "110000010000000000010100101011110100010111111010"; --   -4128748   -5290502
      WHEN  621 => Ti := "110000001000000110010011101011111010100101010011"; --   -4161133   -5265069
      WHEN  622 => Ti := "110000000000001110110000101100000000110101110010"; --   -4193360   -5239438
      WHEN  623 => Ti := "101111111000011001101010101100000111001001010111"; --   -4225430   -5213609
      WHEN  624 => Ti := "101111110000100111000100101100001101100000000000"; --   -4257340   -5187584
      WHEN  625 => Ti := "101111101000110110111101101100010011111001101100"; --   -4289091   -5161364
      WHEN  626 => Ti := "101111100001001001011001101100011010010110011011"; --   -4320679   -5134949
      WHEN  627 => Ti := "101111011001011110010111101100100000110110001010"; --   -4352105   -5108342
      WHEN  628 => Ti := "101111010001110101111000101100100111011000111011"; --   -4383368   -5081541
      WHEN  629 => Ti := "101111001010001111111111101100101101111110101010"; --   -4414465   -5054550
      WHEN  630 => Ti := "101111000010101100101100101100110100100111011000"; --   -4445396   -5027368
      WHEN  631 => Ti := "101110111011001100000000101100111011010011000011"; --   -4476160   -4999997
      WHEN  632 => Ti := "101110110011101101111101101101000010000001101010"; --   -4506755   -4972438
      WHEN  633 => Ti := "101110101100010010100100101101001000110011001101"; --   -4537180   -4944691
      WHEN  634 => Ti := "101110100100111001110101101101001111100111101001"; --   -4567435   -4916759
      WHEN  635 => Ti := "101110011101100011110010101101010110011110111111"; --   -4597518   -4888641
      WHEN  636 => Ti := "101110010110010000011101101101011101011001001101"; --   -4627427   -4860339
      WHEN  637 => Ti := "101110001110111111110101101101100100010110010010"; --   -4657163   -4831854
      WHEN  638 => Ti := "101110000111110001111101101101101011010110001101"; --   -4686723   -4803187
      WHEN  639 => Ti := "101110000000100110110110101101110010011000111100"; --   -4716106   -4774340
      WHEN  640 => Ti := "101101111001011110100000101101111001011110100000"; --   -4745312   -4745312
      WHEN  641 => Ti := "101101110010011000111100101110000000100110110110"; --   -4774340   -4716106
      WHEN  642 => Ti := "101101101011010110001101101110000111110001111101"; --   -4803187   -4686723
      WHEN  643 => Ti := "101101100100010110010010101110001110111111110101"; --   -4831854   -4657163
      WHEN  644 => Ti := "101101011101011001001101101110010110010000011101"; --   -4860339   -4627427
      WHEN  645 => Ti := "101101010110011110111111101110011101100011110010"; --   -4888641   -4597518
      WHEN  646 => Ti := "101101001111100111101001101110100100111001110101"; --   -4916759   -4567435
      WHEN  647 => Ti := "101101001000110011001101101110101100010010100100"; --   -4944691   -4537180
      WHEN  648 => Ti := "101101000010000001101010101110110011101101111101"; --   -4972438   -4506755
      WHEN  649 => Ti := "101100111011010011000011101110111011001100000000"; --   -4999997   -4476160
      WHEN  650 => Ti := "101100110100100111011000101111000010101100101100"; --   -5027368   -4445396
      WHEN  651 => Ti := "101100101101111110101010101111001010001111111111"; --   -5054550   -4414465
      WHEN  652 => Ti := "101100100111011000111011101111010001110101111000"; --   -5081541   -4383368
      WHEN  653 => Ti := "101100100000110110001010101111011001011110010111"; --   -5108342   -4352105
      WHEN  654 => Ti := "101100011010010110011011101111100001001001011001"; --   -5134949   -4320679
      WHEN  655 => Ti := "101100010011111001101100101111101000110110111101"; --   -5161364   -4289091
      WHEN  656 => Ti := "101100001101100000000000101111110000100111000100"; --   -5187584   -4257340
      WHEN  657 => Ti := "101100000111001001010111101111111000011001101010"; --   -5213609   -4225430
      WHEN  658 => Ti := "101100000000110101110010110000000000001110110000"; --   -5239438   -4193360
      WHEN  659 => Ti := "101011111010100101010011110000001000000110010011"; --   -5265069   -4161133
      WHEN  660 => Ti := "101011110100010111111010110000010000000000010100"; --   -5290502   -4128748
      WHEN  661 => Ti := "101011101110001101101000110000010111111100101111"; --   -5315736   -4096209
      WHEN  662 => Ti := "101011101000000110011110110000011111111011100101"; --   -5340770   -4063515
      WHEN  663 => Ti := "101011100010000010011101110000100111111100110100"; --   -5365603   -4030668
      WHEN  664 => Ti := "101011011100000001100111110000110000000000011011"; --   -5390233   -3997669
      WHEN  665 => Ti := "101011010110000011111011110000111000000110011000"; --   -5414661   -3964520
      WHEN  666 => Ti := "101011010000001001011011110001000000001110101010"; --   -5438885   -3931222
      WHEN  667 => Ti := "101011001010010010001000110001001000011001010000"; --   -5462904   -3897776
      WHEN  668 => Ti := "101011000100011110000010110001010000100110001010"; --   -5486718   -3864182
      WHEN  669 => Ti := "101010111110101101001011110001011000110101010100"; --   -5510325   -3830444
      WHEN  670 => Ti := "101010111000111111100100110001100001000110101111"; --   -5533724   -3796561
      WHEN  671 => Ti := "101010110011010101001101110001101001011010011001"; --   -5556915   -3762535
      WHEN  672 => Ti := "101010101101101110000111110001110001110000010000"; --   -5579897   -3728368
      WHEN  673 => Ti := "101010101000001010010011110001111010001000010100"; --   -5602669   -3694060
      WHEN  674 => Ti := "101010100010101001110010110010000010100010100011"; --   -5625230   -3659613
      WHEN  675 => Ti := "101010011101001100100101110010001010111110111100"; --   -5647579   -3625028
      WHEN  676 => Ti := "101010010111110010101101110010010011011101011101"; --   -5669715   -3590307
      WHEN  677 => Ti := "101010010010011100001010110010011011111110000101"; --   -5691638   -3555451
      WHEN  678 => Ti := "101010001101001000111101110010100100100000110011"; --   -5713347   -3520461
      WHEN  679 => Ti := "101010000111111001001000110010101101000101100110"; --   -5734840   -3485338
      WHEN  680 => Ti := "101010000010101100101010110010110101101100011100"; --   -5756118   -3450084
      WHEN  681 => Ti := "101001111101100011100101110010111110010101010100"; --   -5777179   -3414700
      WHEN  682 => Ti := "101001111000011101111010110011000111000000001100"; --   -5798022   -3379188
      WHEN  683 => Ti := "101001110011011011101000110011001111101101000100"; --   -5818648   -3343548
      WHEN  684 => Ti := "101001101110011100110010110011011000011011111001"; --   -5839054   -3307783
      WHEN  685 => Ti := "101001101001100001011000110011100001001100101011"; --   -5859240   -3271893
      WHEN  686 => Ti := "101001100100101001011010110011101001111111011000"; --   -5879206   -3235880
      WHEN  687 => Ti := "101001011111110100111010110011110010110011111111"; --   -5898950   -3199745
      WHEN  688 => Ti := "101001011011000011111000110011111011101010011111"; --   -5918472   -3163489
      WHEN  689 => Ti := "101001010110010110010100110100000100100010110110"; --   -5937772   -3127114
      WHEN  690 => Ti := "101001010001101100010001110100001101011101000010"; --   -5956847   -3090622
      WHEN  691 => Ti := "101001001101000101101101110100010110011001000011"; --   -5975699   -3054013
      WHEN  692 => Ti := "101001001000100010101010110100011111010110110110"; --   -5994326   -3017290
      WHEN  693 => Ti := "101001000100000011001001110100101000010110011100"; --   -6012727   -2980452
      WHEN  694 => Ti := "101000111111100111001011110100110001010111110001"; --   -6030901   -2943503
      WHEN  695 => Ti := "101000111011001110110000110100111010011010110101"; --   -6048848   -2906443
      WHEN  696 => Ti := "101000110110111001111000110101000011011111100111"; --   -6066568   -2869273
      WHEN  697 => Ti := "101000110010101000100100110101001100100110000101"; --   -6084060   -2831995
      WHEN  698 => Ti := "101000101110011010110110110101010101101110001101"; --   -6101322   -2794611
      WHEN  699 => Ti := "101000101010010000101110110101011110110111111111"; --   -6118354   -2757121
      WHEN  700 => Ti := "101000100110001010001011110101101000000011011000"; --   -6135157   -2719528
      WHEN  701 => Ti := "101000100010000111010000110101110001010000011000"; --   -6151728   -2681832
      WHEN  702 => Ti := "101000011110000111111101110101111010011110111101"; --   -6168067   -2644035
      WHEN  703 => Ti := "101000011010001100010001110110000011101111000101"; --   -6184175   -2606139
      WHEN  704 => Ti := "101000010110010100001111110110001101000000110000"; --   -6200049   -2568144
      WHEN  705 => Ti := "101000010010011111110110110110010110010011111011"; --   -6215690   -2530053
      WHEN  706 => Ti := "101000001110101111000110110110011111101000100101"; --   -6231098   -2491867
      WHEN  707 => Ti := "101000001011000010000010110110101000111110101101"; --   -6246270   -2453587
      WHEN  708 => Ti := "101000000111011000101001110110110010010110010010"; --   -6261207   -2415214
      WHEN  709 => Ti := "101000000011110010111011110110111011101111010010"; --   -6275909   -2376750
      WHEN  710 => Ti := "101000000000010000111010110111000101001001101011"; --   -6290374   -2338197
      WHEN  711 => Ti := "100111111100110010100101110111001110100101011100"; --   -6304603   -2299556
      WHEN  712 => Ti := "100111111001010111111110110111011000000010100011"; --   -6318594   -2260829
      WHEN  713 => Ti := "100111110110000001000101110111100001100001000000"; --   -6332347   -2222016
      WHEN  714 => Ti := "100111110010101101111010110111101011000000110000"; --   -6345862   -2183120
      WHEN  715 => Ti := "100111101111011110011110110111110100100001110011"; --   -6359138   -2144141
      WHEN  716 => Ti := "100111101100010010110010110111111110000100000110"; --   -6372174   -2105082
      WHEN  717 => Ti := "100111101001001010110101111000000111100111101001"; --   -6384971   -2065943
      WHEN  718 => Ti := "100111100110000110101001111000010001001100011001"; --   -6397527   -2026727
      WHEN  719 => Ti := "100111100011000110001101111000011010110010010110"; --   -6409843   -1987434
      WHEN  720 => Ti := "100111100000001001100011111000100100011001011101"; --   -6421917   -1948067
      WHEN  721 => Ti := "100111011101010000101011111000101110000001101110"; --   -6433749   -1908626
      WHEN  722 => Ti := "100111011010011011100101111000110111101011000111"; --   -6445339   -1869113
      WHEN  723 => Ti := "100111010111101010010010111001000001010101100110"; --   -6456686   -1829530
      WHEN  724 => Ti := "100111010100111100110010111001001011000001001010"; --   -6467790   -1789878
      WHEN  725 => Ti := "100111010010010011000101111001010100101101110001"; --   -6478651   -1750159
      WHEN  726 => Ti := "100111001111101101001100111001011110011011011010"; --   -6489268   -1710374
      WHEN  727 => Ti := "100111001101001011001000111001101000001010000100"; --   -6499640   -1670524
      WHEN  728 => Ti := "100111001010101100111000111001110001111001101100"; --   -6509768   -1630612
      WHEN  729 => Ti := "100111001000010010011101111001111011101010010010"; --   -6519651   -1590638
      WHEN  730 => Ti := "100111000101111011111000111010000101011011110100"; --   -6529288   -1550604
      WHEN  731 => Ti := "100111000011101001001000111010001111001110010000"; --   -6538680   -1510512
      WHEN  732 => Ti := "100111000001011010001111111010011001000001100101"; --   -6547825   -1470363
      WHEN  733 => Ti := "100110111111001111001100111010100010110101110010"; --   -6556724   -1430158
      WHEN  734 => Ti := "100110111101001000000001111010101100101010110100"; --   -6565375   -1389900
      WHEN  735 => Ti := "100110111011000100101100111010110110100000101010"; --   -6573780   -1349590
      WHEN  736 => Ti := "100110111001000101001111111011000000010111010100"; --   -6581937   -1309228
      WHEN  737 => Ti := "100110110111001001101001111011001010001110101110"; --   -6589847   -1268818
      WHEN  738 => Ti := "100110110101010001111100111011010100000110111001"; --   -6597508   -1228359
      WHEN  739 => Ti := "100110110011011110000111111011011101111111110001"; --   -6604921   -1187855
      WHEN  740 => Ti := "100110110001101110001011111011100111111001010111"; --   -6612085   -1147305
      WHEN  741 => Ti := "100110110000000010001000111011110001110011100111"; --   -6619000   -1106713
      WHEN  742 => Ti := "100110101110011001111110111011111011101110100010"; --   -6625666   -1066078
      WHEN  743 => Ti := "100110101100110101101101111100000101101010000100"; --   -6632083   -1025404
      WHEN  744 => Ti := "100110101011010101010110111100001111100110001101"; --   -6638250    -984691
      WHEN  745 => Ti := "100110101001111000111001111100011001100010111011"; --   -6644167    -943941
      WHEN  746 => Ti := "100110101000100000010110111100100011100000001101"; --   -6649834    -903155
      WHEN  747 => Ti := "100110100111001011101110111100101101011110000000"; --   -6655250    -862336
      WHEN  748 => Ti := "100110100101111011000000111100110111011100010100"; --   -6660416    -821484
      WHEN  749 => Ti := "100110100100101110001101111101000001011011000111"; --   -6665331    -780601
      WHEN  750 => Ti := "100110100011100101010101111101001011011010011000"; --   -6669995    -739688
      WHEN  751 => Ti := "100110100010100000010111111101010101011010000100"; --   -6674409    -698748
      WHEN  752 => Ti := "100110100001011111010110111101011111011010001011"; --   -6678570    -657781
      WHEN  753 => Ti := "100110100000100010001111111101101001011010101010"; --   -6682481    -616790
      WHEN  754 => Ti := "100110011111101001000101111101110011011011100001"; --   -6686139    -575775
      WHEN  755 => Ti := "100110011110110011110110111101111101011100101101"; --   -6689546    -534739
      WHEN  756 => Ti := "100110011110000010100010111110000111011110001101"; --   -6692702    -493683
      WHEN  757 => Ti := "100110011101010101001011111110010001100000000000"; --   -6695605    -452608
      WHEN  758 => Ti := "100110011100101011110000111110011011100010000100"; --   -6698256    -411516
      WHEN  759 => Ti := "100110011100000110010001111110100101100100011000"; --   -6700655    -370408
      WHEN  760 => Ti := "100110011011100100101110111110101111100110111001"; --   -6702802    -329287
      WHEN  761 => Ti := "100110011011000111001000111110111001101001100111"; --   -6704696    -288153
      WHEN  762 => Ti := "100110011010101101011110111111000011101100011111"; --   -6706338    -247009
      WHEN  763 => Ti := "100110011010010111110001111111001101101111100001"; --   -6707727    -205855
      WHEN  764 => Ti := "100110011010000110000000111111010111110010101011"; --   -6708864    -164693
      WHEN  765 => Ti := "100110011001111000001100111111100001110101111011"; --   -6709748    -123525
      WHEN  766 => Ti := "100110011001101110010100111111101011111001010000"; --   -6710380     -82352
      WHEN  767 => Ti := "100110011001101000011001111111110101111100100111"; --   -6710759     -41177
      WHEN  768 => Ti := "100110011001100110011011000000000000000000000000"; --   -6710885         +0
      WHEN  769 => Ti := "100110011001101000011001000000001010000011011001"; --   -6710759     +41177
      WHEN  770 => Ti := "100110011001101110010100000000010100000110110000"; --   -6710380     +82352
      WHEN  771 => Ti := "100110011001111000001100000000011110001010000101"; --   -6709748    +123525
      WHEN  772 => Ti := "100110011010000110000000000000101000001101010101"; --   -6708864    +164693
      WHEN  773 => Ti := "100110011010010111110001000000110010010000011111"; --   -6707727    +205855
      WHEN  774 => Ti := "100110011010101101011110000000111100010011100001"; --   -6706338    +247009
      WHEN  775 => Ti := "100110011011000111001000000001000110010110011001"; --   -6704696    +288153
      WHEN  776 => Ti := "100110011011100100101110000001010000011001000111"; --   -6702802    +329287
      WHEN  777 => Ti := "100110011100000110010001000001011010011011101000"; --   -6700655    +370408
      WHEN  778 => Ti := "100110011100101011110000000001100100011101111100"; --   -6698256    +411516
      WHEN  779 => Ti := "100110011101010101001011000001101110100000000000"; --   -6695605    +452608
      WHEN  780 => Ti := "100110011110000010100010000001111000100001110011"; --   -6692702    +493683
      WHEN  781 => Ti := "100110011110110011110110000010000010100011010011"; --   -6689546    +534739
      WHEN  782 => Ti := "100110011111101001000101000010001100100100011111"; --   -6686139    +575775
      WHEN  783 => Ti := "100110100000100010001111000010010110100101010110"; --   -6682481    +616790
      WHEN  784 => Ti := "100110100001011111010110000010100000100101110101"; --   -6678570    +657781
      WHEN  785 => Ti := "100110100010100000010111000010101010100101111100"; --   -6674409    +698748
      WHEN  786 => Ti := "100110100011100101010101000010110100100101101000"; --   -6669995    +739688
      WHEN  787 => Ti := "100110100100101110001101000010111110100100111001"; --   -6665331    +780601
      WHEN  788 => Ti := "100110100101111011000000000011001000100011101100"; --   -6660416    +821484
      WHEN  789 => Ti := "100110100111001011101110000011010010100010000000"; --   -6655250    +862336
      WHEN  790 => Ti := "100110101000100000010110000011011100011111110011"; --   -6649834    +903155
      WHEN  791 => Ti := "100110101001111000111001000011100110011101000101"; --   -6644167    +943941
      WHEN  792 => Ti := "100110101011010101010110000011110000011001110011"; --   -6638250    +984691
      WHEN  793 => Ti := "100110101100110101101101000011111010010101111100"; --   -6632083   +1025404
      WHEN  794 => Ti := "100110101110011001111110000100000100010001011110"; --   -6625666   +1066078
      WHEN  795 => Ti := "100110110000000010001000000100001110001100011001"; --   -6619000   +1106713
      WHEN  796 => Ti := "100110110001101110001011000100011000000110101001"; --   -6612085   +1147305
      WHEN  797 => Ti := "100110110011011110000111000100100010000000001111"; --   -6604921   +1187855
      WHEN  798 => Ti := "100110110101010001111100000100101011111001000111"; --   -6597508   +1228359
      WHEN  799 => Ti := "100110110111001001101001000100110101110001010010"; --   -6589847   +1268818
      WHEN  800 => Ti := "100110111001000101001111000100111111101000101100"; --   -6581937   +1309228
      WHEN  801 => Ti := "100110111011000100101100000101001001011111010110"; --   -6573780   +1349590
      WHEN  802 => Ti := "100110111101001000000001000101010011010101001100"; --   -6565375   +1389900
      WHEN  803 => Ti := "100110111111001111001100000101011101001010001110"; --   -6556724   +1430158
      WHEN  804 => Ti := "100111000001011010001111000101100110111110011011"; --   -6547825   +1470363
      WHEN  805 => Ti := "100111000011101001001000000101110000110001110000"; --   -6538680   +1510512
      WHEN  806 => Ti := "100111000101111011111000000101111010100100001100"; --   -6529288   +1550604
      WHEN  807 => Ti := "100111001000010010011101000110000100010101101110"; --   -6519651   +1590638
      WHEN  808 => Ti := "100111001010101100111000000110001110000110010100"; --   -6509768   +1630612
      WHEN  809 => Ti := "100111001101001011001000000110010111110101111100"; --   -6499640   +1670524
      WHEN  810 => Ti := "100111001111101101001100000110100001100100100110"; --   -6489268   +1710374
      WHEN  811 => Ti := "100111010010010011000101000110101011010010001111"; --   -6478651   +1750159
      WHEN  812 => Ti := "100111010100111100110010000110110100111110110110"; --   -6467790   +1789878
      WHEN  813 => Ti := "100111010111101010010010000110111110101010011010"; --   -6456686   +1829530
      WHEN  814 => Ti := "100111011010011011100101000111001000010100111001"; --   -6445339   +1869113
      WHEN  815 => Ti := "100111011101010000101011000111010001111110010010"; --   -6433749   +1908626
      WHEN  816 => Ti := "100111100000001001100011000111011011100110100011"; --   -6421917   +1948067
      WHEN  817 => Ti := "100111100011000110001101000111100101001101101010"; --   -6409843   +1987434
      WHEN  818 => Ti := "100111100110000110101001000111101110110011100111"; --   -6397527   +2026727
      WHEN  819 => Ti := "100111101001001010110101000111111000011000010111"; --   -6384971   +2065943
      WHEN  820 => Ti := "100111101100010010110010001000000001111011111010"; --   -6372174   +2105082
      WHEN  821 => Ti := "100111101111011110011110001000001011011110001101"; --   -6359138   +2144141
      WHEN  822 => Ti := "100111110010101101111010001000010100111111010000"; --   -6345862   +2183120
      WHEN  823 => Ti := "100111110110000001000101001000011110011111000000"; --   -6332347   +2222016
      WHEN  824 => Ti := "100111111001010111111110001000100111111101011101"; --   -6318594   +2260829
      WHEN  825 => Ti := "100111111100110010100101001000110001011010100100"; --   -6304603   +2299556
      WHEN  826 => Ti := "101000000000010000111010001000111010110110010101"; --   -6290374   +2338197
      WHEN  827 => Ti := "101000000011110010111011001001000100010000101110"; --   -6275909   +2376750
      WHEN  828 => Ti := "101000000111011000101001001001001101101001101110"; --   -6261207   +2415214
      WHEN  829 => Ti := "101000001011000010000010001001010111000001010011"; --   -6246270   +2453587
      WHEN  830 => Ti := "101000001110101111000110001001100000010111011011"; --   -6231098   +2491867
      WHEN  831 => Ti := "101000010010011111110110001001101001101100000101"; --   -6215690   +2530053
      WHEN  832 => Ti := "101000010110010100001111001001110010111111010000"; --   -6200049   +2568144
      WHEN  833 => Ti := "101000011010001100010001001001111100010000111011"; --   -6184175   +2606139
      WHEN  834 => Ti := "101000011110000111111101001010000101100001000011"; --   -6168067   +2644035
      WHEN  835 => Ti := "101000100010000111010000001010001110101111101000"; --   -6151728   +2681832
      WHEN  836 => Ti := "101000100110001010001011001010010111111100101000"; --   -6135157   +2719528
      WHEN  837 => Ti := "101000101010010000101110001010100001001000000001"; --   -6118354   +2757121
      WHEN  838 => Ti := "101000101110011010110110001010101010010001110011"; --   -6101322   +2794611
      WHEN  839 => Ti := "101000110010101000100100001010110011011001111011"; --   -6084060   +2831995
      WHEN  840 => Ti := "101000110110111001111000001010111100100000011001"; --   -6066568   +2869273
      WHEN  841 => Ti := "101000111011001110110000001011000101100101001011"; --   -6048848   +2906443
      WHEN  842 => Ti := "101000111111100111001011001011001110101000001111"; --   -6030901   +2943503
      WHEN  843 => Ti := "101001000100000011001001001011010111101001100100"; --   -6012727   +2980452
      WHEN  844 => Ti := "101001001000100010101010001011100000101001001010"; --   -5994326   +3017290
      WHEN  845 => Ti := "101001001101000101101101001011101001100110111101"; --   -5975699   +3054013
      WHEN  846 => Ti := "101001010001101100010001001011110010100010111110"; --   -5956847   +3090622
      WHEN  847 => Ti := "101001010110010110010100001011111011011101001010"; --   -5937772   +3127114
      WHEN  848 => Ti := "101001011011000011111000001100000100010101100001"; --   -5918472   +3163489
      WHEN  849 => Ti := "101001011111110100111010001100001101001100000001"; --   -5898950   +3199745
      WHEN  850 => Ti := "101001100100101001011010001100010110000000101000"; --   -5879206   +3235880
      WHEN  851 => Ti := "101001101001100001011000001100011110110011010101"; --   -5859240   +3271893
      WHEN  852 => Ti := "101001101110011100110010001100100111100100000111"; --   -5839054   +3307783
      WHEN  853 => Ti := "101001110011011011101000001100110000010010111100"; --   -5818648   +3343548
      WHEN  854 => Ti := "101001111000011101111010001100111000111111110100"; --   -5798022   +3379188
      WHEN  855 => Ti := "101001111101100011100101001101000001101010101100"; --   -5777179   +3414700
      WHEN  856 => Ti := "101010000010101100101010001101001010010011100100"; --   -5756118   +3450084
      WHEN  857 => Ti := "101010000111111001001000001101010010111010011010"; --   -5734840   +3485338
      WHEN  858 => Ti := "101010001101001000111101001101011011011111001101"; --   -5713347   +3520461
      WHEN  859 => Ti := "101010010010011100001010001101100100000001111011"; --   -5691638   +3555451
      WHEN  860 => Ti := "101010010111110010101101001101101100100010100011"; --   -5669715   +3590307
      WHEN  861 => Ti := "101010011101001100100101001101110101000001000100"; --   -5647579   +3625028
      WHEN  862 => Ti := "101010100010101001110010001101111101011101011101"; --   -5625230   +3659613
      WHEN  863 => Ti := "101010101000001010010011001110000101110111101100"; --   -5602669   +3694060
      WHEN  864 => Ti := "101010101101101110000111001110001110001111110000"; --   -5579897   +3728368
      WHEN  865 => Ti := "101010110011010101001101001110010110100101100111"; --   -5556915   +3762535
      WHEN  866 => Ti := "101010111000111111100100001110011110111001010001"; --   -5533724   +3796561
      WHEN  867 => Ti := "101010111110101101001011001110100111001010101100"; --   -5510325   +3830444
      WHEN  868 => Ti := "101011000100011110000010001110101111011001110110"; --   -5486718   +3864182
      WHEN  869 => Ti := "101011001010010010001000001110110111100110110000"; --   -5462904   +3897776
      WHEN  870 => Ti := "101011010000001001011011001110111111110001010110"; --   -5438885   +3931222
      WHEN  871 => Ti := "101011010110000011111011001111000111111001101000"; --   -5414661   +3964520
      WHEN  872 => Ti := "101011011100000001100111001111001111111111100101"; --   -5390233   +3997669
      WHEN  873 => Ti := "101011100010000010011101001111011000000011001100"; --   -5365603   +4030668
      WHEN  874 => Ti := "101011101000000110011110001111100000000100011011"; --   -5340770   +4063515
      WHEN  875 => Ti := "101011101110001101101000001111101000000011010001"; --   -5315736   +4096209
      WHEN  876 => Ti := "101011110100010111111010001111101111111111101100"; --   -5290502   +4128748
      WHEN  877 => Ti := "101011111010100101010011001111110111111001101101"; --   -5265069   +4161133
      WHEN  878 => Ti := "101100000000110101110010001111111111110001010000"; --   -5239438   +4193360
      WHEN  879 => Ti := "101100000111001001010111010000000111100110010110"; --   -5213609   +4225430
      WHEN  880 => Ti := "101100001101100000000000010000001111011000111100"; --   -5187584   +4257340
      WHEN  881 => Ti := "101100010011111001101100010000010111001001000011"; --   -5161364   +4289091
      WHEN  882 => Ti := "101100011010010110011011010000011110110110100111"; --   -5134949   +4320679
      WHEN  883 => Ti := "101100100000110110001010010000100110100001101001"; --   -5108342   +4352105
      WHEN  884 => Ti := "101100100111011000111011010000101110001010001000"; --   -5081541   +4383368
      WHEN  885 => Ti := "101100101101111110101010010000110101110000000001"; --   -5054550   +4414465
      WHEN  886 => Ti := "101100110100100111011000010000111101010011010100"; --   -5027368   +4445396
      WHEN  887 => Ti := "101100111011010011000011010001000100110100000000"; --   -4999997   +4476160
      WHEN  888 => Ti := "101101000010000001101010010001001100010010000011"; --   -4972438   +4506755
      WHEN  889 => Ti := "101101001000110011001101010001010011101101011100"; --   -4944691   +4537180
      WHEN  890 => Ti := "101101001111100111101001010001011011000110001011"; --   -4916759   +4567435
      WHEN  891 => Ti := "101101010110011110111111010001100010011100001110"; --   -4888641   +4597518
      WHEN  892 => Ti := "101101011101011001001101010001101001101111100011"; --   -4860339   +4627427
      WHEN  893 => Ti := "101101100100010110010010010001110001000000001011"; --   -4831854   +4657163
      WHEN  894 => Ti := "101101101011010110001101010001111000001110000011"; --   -4803187   +4686723
      WHEN  895 => Ti := "101101110010011000111100010001111111011001001010"; --   -4774340   +4716106
      WHEN  896 => Ti := "101101111001011110100000010010000110100001100000"; --   -4745312   +4745312
      WHEN  897 => Ti := "101110000000100110110110010010001101100111000100"; --   -4716106   +4774340
      WHEN  898 => Ti := "101110000111110001111101010010010100101001110011"; --   -4686723   +4803187
      WHEN  899 => Ti := "101110001110111111110101010010011011101001101110"; --   -4657163   +4831854
      WHEN  900 => Ti := "101110010110010000011101010010100010100110110011"; --   -4627427   +4860339
      WHEN  901 => Ti := "101110011101100011110010010010101001100001000001"; --   -4597518   +4888641
      WHEN  902 => Ti := "101110100100111001110101010010110000011000010111"; --   -4567435   +4916759
      WHEN  903 => Ti := "101110101100010010100100010010110111001100110011"; --   -4537180   +4944691
      WHEN  904 => Ti := "101110110011101101111101010010111101111110010110"; --   -4506755   +4972438
      WHEN  905 => Ti := "101110111011001100000000010011000100101100111101"; --   -4476160   +4999997
      WHEN  906 => Ti := "101111000010101100101100010011001011011000101000"; --   -4445396   +5027368
      WHEN  907 => Ti := "101111001010001111111111010011010010000001010110"; --   -4414465   +5054550
      WHEN  908 => Ti := "101111010001110101111000010011011000100111000101"; --   -4383368   +5081541
      WHEN  909 => Ti := "101111011001011110010111010011011111001001110110"; --   -4352105   +5108342
      WHEN  910 => Ti := "101111100001001001011001010011100101101001100101"; --   -4320679   +5134949
      WHEN  911 => Ti := "101111101000110110111101010011101100000110010100"; --   -4289091   +5161364
      WHEN  912 => Ti := "101111110000100111000100010011110010100000000000"; --   -4257340   +5187584
      WHEN  913 => Ti := "101111111000011001101010010011111000110110101001"; --   -4225430   +5213609
      WHEN  914 => Ti := "110000000000001110110000010011111111001010001110"; --   -4193360   +5239438
      WHEN  915 => Ti := "110000001000000110010011010100000101011010101101"; --   -4161133   +5265069
      WHEN  916 => Ti := "110000010000000000010100010100001011101000000110"; --   -4128748   +5290502
      WHEN  917 => Ti := "110000010111111100101111010100010001110010011000"; --   -4096209   +5315736
      WHEN  918 => Ti := "110000011111111011100101010100010111111001100010"; --   -4063515   +5340770
      WHEN  919 => Ti := "110000100111111100110100010100011101111101100011"; --   -4030668   +5365603
      WHEN  920 => Ti := "110000110000000000011011010100100011111110011001"; --   -3997669   +5390233
      WHEN  921 => Ti := "110000111000000110011000010100101001111100000101"; --   -3964520   +5414661
      WHEN  922 => Ti := "110001000000001110101010010100101111110110100101"; --   -3931222   +5438885
      WHEN  923 => Ti := "110001001000011001010000010100110101101101111000"; --   -3897776   +5462904
      WHEN  924 => Ti := "110001010000100110001010010100111011100001111110"; --   -3864182   +5486718
      WHEN  925 => Ti := "110001011000110101010100010101000001010010110101"; --   -3830444   +5510325
      WHEN  926 => Ti := "110001100001000110101111010101000111000000011100"; --   -3796561   +5533724
      WHEN  927 => Ti := "110001101001011010011001010101001100101010110011"; --   -3762535   +5556915
      WHEN  928 => Ti := "110001110001110000010000010101010010010001111001"; --   -3728368   +5579897
      WHEN  929 => Ti := "110001111010001000010100010101010111110101101101"; --   -3694060   +5602669
      WHEN  930 => Ti := "110010000010100010100011010101011101010110001110"; --   -3659613   +5625230
      WHEN  931 => Ti := "110010001010111110111100010101100010110011011011"; --   -3625028   +5647579
      WHEN  932 => Ti := "110010010011011101011101010101101000001101010011"; --   -3590307   +5669715
      WHEN  933 => Ti := "110010011011111110000101010101101101100011110110"; --   -3555451   +5691638
      WHEN  934 => Ti := "110010100100100000110011010101110010110111000011"; --   -3520461   +5713347
      WHEN  935 => Ti := "110010101101000101100110010101111000000110111000"; --   -3485338   +5734840
      WHEN  936 => Ti := "110010110101101100011100010101111101010011010110"; --   -3450084   +5756118
      WHEN  937 => Ti := "110010111110010101010100010110000010011100011011"; --   -3414700   +5777179
      WHEN  938 => Ti := "110011000111000000001100010110000111100010000110"; --   -3379188   +5798022
      WHEN  939 => Ti := "110011001111101101000100010110001100100100011000"; --   -3343548   +5818648
      WHEN  940 => Ti := "110011011000011011111001010110010001100011001110"; --   -3307783   +5839054
      WHEN  941 => Ti := "110011100001001100101011010110010110011110101000"; --   -3271893   +5859240
      WHEN  942 => Ti := "110011101001111111011000010110011011010110100110"; --   -3235880   +5879206
      WHEN  943 => Ti := "110011110010110011111111010110100000001011000110"; --   -3199745   +5898950
      WHEN  944 => Ti := "110011111011101010011111010110100100111100001000"; --   -3163489   +5918472
      WHEN  945 => Ti := "110100000100100010110110010110101001101001101100"; --   -3127114   +5937772
      WHEN  946 => Ti := "110100001101011101000010010110101110010011101111"; --   -3090622   +5956847
      WHEN  947 => Ti := "110100010110011001000011010110110010111010010011"; --   -3054013   +5975699
      WHEN  948 => Ti := "110100011111010110110110010110110111011101010110"; --   -3017290   +5994326
      WHEN  949 => Ti := "110100101000010110011100010110111011111100110111"; --   -2980452   +6012727
      WHEN  950 => Ti := "110100110001010111110001010111000000011000110101"; --   -2943503   +6030901
      WHEN  951 => Ti := "110100111010011010110101010111000100110001010000"; --   -2906443   +6048848
      WHEN  952 => Ti := "110101000011011111100111010111001001000110001000"; --   -2869273   +6066568
      WHEN  953 => Ti := "110101001100100110000101010111001101010111011100"; --   -2831995   +6084060
      WHEN  954 => Ti := "110101010101101110001101010111010001100101001010"; --   -2794611   +6101322
      WHEN  955 => Ti := "110101011110110111111111010111010101101111010010"; --   -2757121   +6118354
      WHEN  956 => Ti := "110101101000000011011000010111011001110101110101"; --   -2719528   +6135157
      WHEN  957 => Ti := "110101110001010000011000010111011101111000110000"; --   -2681832   +6151728
      WHEN  958 => Ti := "110101111010011110111101010111100001111000000011"; --   -2644035   +6168067
      WHEN  959 => Ti := "110110000011101111000101010111100101110011101111"; --   -2606139   +6184175
      WHEN  960 => Ti := "110110001101000000110000010111101001101011110001"; --   -2568144   +6200049
      WHEN  961 => Ti := "110110010110010011111011010111101101100000001010"; --   -2530053   +6215690
      WHEN  962 => Ti := "110110011111101000100101010111110001010000111010"; --   -2491867   +6231098
      WHEN  963 => Ti := "110110101000111110101101010111110100111101111110"; --   -2453587   +6246270
      WHEN  964 => Ti := "110110110010010110010010010111111000100111010111"; --   -2415214   +6261207
      WHEN  965 => Ti := "110110111011101111010010010111111100001101000101"; --   -2376750   +6275909
      WHEN  966 => Ti := "110111000101001001101011010111111111101111000110"; --   -2338197   +6290374
      WHEN  967 => Ti := "110111001110100101011100011000000011001101011011"; --   -2299556   +6304603
      WHEN  968 => Ti := "110111011000000010100011011000000110101000000010"; --   -2260829   +6318594
      WHEN  969 => Ti := "110111100001100001000000011000001001111110111011"; --   -2222016   +6332347
      WHEN  970 => Ti := "110111101011000000110000011000001101010010000110"; --   -2183120   +6345862
      WHEN  971 => Ti := "110111110100100001110011011000010000100001100010"; --   -2144141   +6359138
      WHEN  972 => Ti := "110111111110000100000110011000010011101101001110"; --   -2105082   +6372174
      WHEN  973 => Ti := "111000000111100111101001011000010110110101001011"; --   -2065943   +6384971
      WHEN  974 => Ti := "111000010001001100011001011000011001111001010111"; --   -2026727   +6397527
      WHEN  975 => Ti := "111000011010110010010110011000011100111001110011"; --   -1987434   +6409843
      WHEN  976 => Ti := "111000100100011001011101011000011111110110011101"; --   -1948067   +6421917
      WHEN  977 => Ti := "111000101110000001101110011000100010101111010101"; --   -1908626   +6433749
      WHEN  978 => Ti := "111000110111101011000111011000100101100100011011"; --   -1869113   +6445339
      WHEN  979 => Ti := "111001000001010101100110011000101000010101101110"; --   -1829530   +6456686
      WHEN  980 => Ti := "111001001011000001001010011000101011000011001110"; --   -1789878   +6467790
      WHEN  981 => Ti := "111001010100101101110001011000101101101100111011"; --   -1750159   +6478651
      WHEN  982 => Ti := "111001011110011011011010011000110000010010110100"; --   -1710374   +6489268
      WHEN  983 => Ti := "111001101000001010000100011000110010110100111000"; --   -1670524   +6499640
      WHEN  984 => Ti := "111001110001111001101100011000110101010011001000"; --   -1630612   +6509768
      WHEN  985 => Ti := "111001111011101010010010011000110111101101100011"; --   -1590638   +6519651
      WHEN  986 => Ti := "111010000101011011110100011000111010000100001000"; --   -1550604   +6529288
      WHEN  987 => Ti := "111010001111001110010000011000111100010110111000"; --   -1510512   +6538680
      WHEN  988 => Ti := "111010011001000001100101011000111110100101110001"; --   -1470363   +6547825
      WHEN  989 => Ti := "111010100010110101110010011001000000110000110100"; --   -1430158   +6556724
      WHEN  990 => Ti := "111010101100101010110100011001000010110111111111"; --   -1389900   +6565375
      WHEN  991 => Ti := "111010110110100000101010011001000100111011010100"; --   -1349590   +6573780
      WHEN  992 => Ti := "111011000000010111010100011001000110111010110001"; --   -1309228   +6581937
      WHEN  993 => Ti := "111011001010001110101110011001001000110110010111"; --   -1268818   +6589847
      WHEN  994 => Ti := "111011010100000110111001011001001010101110000100"; --   -1228359   +6597508
      WHEN  995 => Ti := "111011011101111111110001011001001100100001111001"; --   -1187855   +6604921
      WHEN  996 => Ti := "111011100111111001010111011001001110010001110101"; --   -1147305   +6612085
      WHEN  997 => Ti := "111011110001110011100111011001001111111101111000"; --   -1106713   +6619000
      WHEN  998 => Ti := "111011111011101110100010011001010001100110000010"; --   -1066078   +6625666
      WHEN  999 => Ti := "111100000101101010000100011001010011001010010011"; --   -1025404   +6632083
      WHEN 1000 => Ti := "111100001111100110001101011001010100101010101010"; --    -984691   +6638250
      WHEN 1001 => Ti := "111100011001100010111011011001010110000111000111"; --    -943941   +6644167
      WHEN 1002 => Ti := "111100100011100000001101011001010111011111101010"; --    -903155   +6649834
      WHEN 1003 => Ti := "111100101101011110000000011001011000110100010010"; --    -862336   +6655250
      WHEN 1004 => Ti := "111100110111011100010100011001011010000101000000"; --    -821484   +6660416
      WHEN 1005 => Ti := "111101000001011011000111011001011011010001110011"; --    -780601   +6665331
      WHEN 1006 => Ti := "111101001011011010011000011001011100011010101011"; --    -739688   +6669995
      WHEN 1007 => Ti := "111101010101011010000100011001011101011111101001"; --    -698748   +6674409
      WHEN 1008 => Ti := "111101011111011010001011011001011110100000101010"; --    -657781   +6678570
      WHEN 1009 => Ti := "111101101001011010101010011001011111011101110001"; --    -616790   +6682481
      WHEN 1010 => Ti := "111101110011011011100001011001100000010110111011"; --    -575775   +6686139
      WHEN 1011 => Ti := "111101111101011100101101011001100001001100001010"; --    -534739   +6689546
      WHEN 1012 => Ti := "111110000111011110001101011001100001111101011110"; --    -493683   +6692702
      WHEN 1013 => Ti := "111110010001100000000000011001100010101010110101"; --    -452608   +6695605
      WHEN 1014 => Ti := "111110011011100010000100011001100011010100010000"; --    -411516   +6698256
      WHEN 1015 => Ti := "111110100101100100011000011001100011111001101111"; --    -370408   +6700655
      WHEN 1016 => Ti := "111110101111100110111001011001100100011011010010"; --    -329287   +6702802
      WHEN 1017 => Ti := "111110111001101001100111011001100100111000111000"; --    -288153   +6704696
      WHEN 1018 => Ti := "111111000011101100011111011001100101010010100010"; --    -247009   +6706338
      WHEN 1019 => Ti := "111111001101101111100001011001100101101000001111"; --    -205855   +6707727
      WHEN 1020 => Ti := "111111010111110010101011011001100101111010000000"; --    -164693   +6708864
      WHEN 1021 => Ti := "111111100001110101111011011001100110000111110100"; --    -123525   +6709748
      WHEN 1022 => Ti := "111111101011111001010000011001100110010001101100"; --     -82352   +6710380
      WHEN 1023 => Ti := "111111110101111100100111011001100110010111100111"; --     -41177   +6710759
      WHEN 1024 => Ti := "000000000000000000000000011001100110011001100101"; --         +0   +6710885
      WHEN 1025 => Ti := "000000001010000011011001011001100110010111100111"; --     +41177   +6710759
      WHEN 1026 => Ti := "000000010100000110110000011001100110010001101100"; --     +82352   +6710380
      WHEN 1027 => Ti := "000000011110001010000101011001100110000111110100"; --    +123525   +6709748
      WHEN 1028 => Ti := "000000101000001101010101011001100101111010000000"; --    +164693   +6708864
      WHEN 1029 => Ti := "000000110010010000011111011001100101101000001111"; --    +205855   +6707727
      WHEN 1030 => Ti := "000000111100010011100001011001100101010010100010"; --    +247009   +6706338
      WHEN 1031 => Ti := "000001000110010110011001011001100100111000111000"; --    +288153   +6704696
      WHEN 1032 => Ti := "000001010000011001000111011001100100011011010010"; --    +329287   +6702802
      WHEN 1033 => Ti := "000001011010011011101000011001100011111001101111"; --    +370408   +6700655
      WHEN 1034 => Ti := "000001100100011101111100011001100011010100010000"; --    +411516   +6698256
      WHEN 1035 => Ti := "000001101110100000000000011001100010101010110101"; --    +452608   +6695605
      WHEN 1036 => Ti := "000001111000100001110011011001100001111101011110"; --    +493683   +6692702
      WHEN 1037 => Ti := "000010000010100011010011011001100001001100001010"; --    +534739   +6689546
      WHEN 1038 => Ti := "000010001100100100011111011001100000010110111011"; --    +575775   +6686139
      WHEN 1039 => Ti := "000010010110100101010110011001011111011101110001"; --    +616790   +6682481
      WHEN 1040 => Ti := "000010100000100101110101011001011110100000101010"; --    +657781   +6678570
      WHEN 1041 => Ti := "000010101010100101111100011001011101011111101001"; --    +698748   +6674409
      WHEN 1042 => Ti := "000010110100100101101000011001011100011010101011"; --    +739688   +6669995
      WHEN 1043 => Ti := "000010111110100100111001011001011011010001110011"; --    +780601   +6665331
      WHEN 1044 => Ti := "000011001000100011101100011001011010000101000000"; --    +821484   +6660416
      WHEN 1045 => Ti := "000011010010100010000000011001011000110100010010"; --    +862336   +6655250
      WHEN 1046 => Ti := "000011011100011111110011011001010111011111101010"; --    +903155   +6649834
      WHEN 1047 => Ti := "000011100110011101000101011001010110000111000111"; --    +943941   +6644167
      WHEN 1048 => Ti := "000011110000011001110011011001010100101010101010"; --    +984691   +6638250
      WHEN 1049 => Ti := "000011111010010101111100011001010011001010010011"; --   +1025404   +6632083
      WHEN 1050 => Ti := "000100000100010001011110011001010001100110000010"; --   +1066078   +6625666
      WHEN 1051 => Ti := "000100001110001100011001011001001111111101111000"; --   +1106713   +6619000
      WHEN 1052 => Ti := "000100011000000110101001011001001110010001110101"; --   +1147305   +6612085
      WHEN 1053 => Ti := "000100100010000000001111011001001100100001111001"; --   +1187855   +6604921
      WHEN 1054 => Ti := "000100101011111001000111011001001010101110000100"; --   +1228359   +6597508
      WHEN 1055 => Ti := "000100110101110001010010011001001000110110010111"; --   +1268818   +6589847
      WHEN 1056 => Ti := "000100111111101000101100011001000110111010110001"; --   +1309228   +6581937
      WHEN 1057 => Ti := "000101001001011111010110011001000100111011010100"; --   +1349590   +6573780
      WHEN 1058 => Ti := "000101010011010101001100011001000010110111111111"; --   +1389900   +6565375
      WHEN 1059 => Ti := "000101011101001010001110011001000000110000110100"; --   +1430158   +6556724
      WHEN 1060 => Ti := "000101100110111110011011011000111110100101110001"; --   +1470363   +6547825
      WHEN 1061 => Ti := "000101110000110001110000011000111100010110111000"; --   +1510512   +6538680
      WHEN 1062 => Ti := "000101111010100100001100011000111010000100001000"; --   +1550604   +6529288
      WHEN 1063 => Ti := "000110000100010101101110011000110111101101100011"; --   +1590638   +6519651
      WHEN 1064 => Ti := "000110001110000110010100011000110101010011001000"; --   +1630612   +6509768
      WHEN 1065 => Ti := "000110010111110101111100011000110010110100111000"; --   +1670524   +6499640
      WHEN 1066 => Ti := "000110100001100100100110011000110000010010110100"; --   +1710374   +6489268
      WHEN 1067 => Ti := "000110101011010010001111011000101101101100111011"; --   +1750159   +6478651
      WHEN 1068 => Ti := "000110110100111110110110011000101011000011001110"; --   +1789878   +6467790
      WHEN 1069 => Ti := "000110111110101010011010011000101000010101101110"; --   +1829530   +6456686
      WHEN 1070 => Ti := "000111001000010100111001011000100101100100011011"; --   +1869113   +6445339
      WHEN 1071 => Ti := "000111010001111110010010011000100010101111010101"; --   +1908626   +6433749
      WHEN 1072 => Ti := "000111011011100110100011011000011111110110011101"; --   +1948067   +6421917
      WHEN 1073 => Ti := "000111100101001101101010011000011100111001110011"; --   +1987434   +6409843
      WHEN 1074 => Ti := "000111101110110011100111011000011001111001010111"; --   +2026727   +6397527
      WHEN 1075 => Ti := "000111111000011000010111011000010110110101001011"; --   +2065943   +6384971
      WHEN 1076 => Ti := "001000000001111011111010011000010011101101001110"; --   +2105082   +6372174
      WHEN 1077 => Ti := "001000001011011110001101011000010000100001100010"; --   +2144141   +6359138
      WHEN 1078 => Ti := "001000010100111111010000011000001101010010000110"; --   +2183120   +6345862
      WHEN 1079 => Ti := "001000011110011111000000011000001001111110111011"; --   +2222016   +6332347
      WHEN 1080 => Ti := "001000100111111101011101011000000110101000000010"; --   +2260829   +6318594
      WHEN 1081 => Ti := "001000110001011010100100011000000011001101011011"; --   +2299556   +6304603
      WHEN 1082 => Ti := "001000111010110110010101010111111111101111000110"; --   +2338197   +6290374
      WHEN 1083 => Ti := "001001000100010000101110010111111100001101000101"; --   +2376750   +6275909
      WHEN 1084 => Ti := "001001001101101001101110010111111000100111010111"; --   +2415214   +6261207
      WHEN 1085 => Ti := "001001010111000001010011010111110100111101111110"; --   +2453587   +6246270
      WHEN 1086 => Ti := "001001100000010111011011010111110001010000111010"; --   +2491867   +6231098
      WHEN 1087 => Ti := "001001101001101100000101010111101101100000001010"; --   +2530053   +6215690
      WHEN 1088 => Ti := "001001110010111111010000010111101001101011110001"; --   +2568144   +6200049
      WHEN 1089 => Ti := "001001111100010000111011010111100101110011101111"; --   +2606139   +6184175
      WHEN 1090 => Ti := "001010000101100001000011010111100001111000000011"; --   +2644035   +6168067
      WHEN 1091 => Ti := "001010001110101111101000010111011101111000110000"; --   +2681832   +6151728
      WHEN 1092 => Ti := "001010010111111100101000010111011001110101110101"; --   +2719528   +6135157
      WHEN 1093 => Ti := "001010100001001000000001010111010101101111010010"; --   +2757121   +6118354
      WHEN 1094 => Ti := "001010101010010001110011010111010001100101001010"; --   +2794611   +6101322
      WHEN 1095 => Ti := "001010110011011001111011010111001101010111011100"; --   +2831995   +6084060
      WHEN 1096 => Ti := "001010111100100000011001010111001001000110001000"; --   +2869273   +6066568
      WHEN 1097 => Ti := "001011000101100101001011010111000100110001010000"; --   +2906443   +6048848
      WHEN 1098 => Ti := "001011001110101000001111010111000000011000110101"; --   +2943503   +6030901
      WHEN 1099 => Ti := "001011010111101001100100010110111011111100110111"; --   +2980452   +6012727
      WHEN 1100 => Ti := "001011100000101001001010010110110111011101010110"; --   +3017290   +5994326
      WHEN 1101 => Ti := "001011101001100110111101010110110010111010010011"; --   +3054013   +5975699
      WHEN 1102 => Ti := "001011110010100010111110010110101110010011101111"; --   +3090622   +5956847
      WHEN 1103 => Ti := "001011111011011101001010010110101001101001101100"; --   +3127114   +5937772
      WHEN 1104 => Ti := "001100000100010101100001010110100100111100001000"; --   +3163489   +5918472
      WHEN 1105 => Ti := "001100001101001100000001010110100000001011000110"; --   +3199745   +5898950
      WHEN 1106 => Ti := "001100010110000000101000010110011011010110100110"; --   +3235880   +5879206
      WHEN 1107 => Ti := "001100011110110011010101010110010110011110101000"; --   +3271893   +5859240
      WHEN 1108 => Ti := "001100100111100100000111010110010001100011001110"; --   +3307783   +5839054
      WHEN 1109 => Ti := "001100110000010010111100010110001100100100011000"; --   +3343548   +5818648
      WHEN 1110 => Ti := "001100111000111111110100010110000111100010000110"; --   +3379188   +5798022
      WHEN 1111 => Ti := "001101000001101010101100010110000010011100011011"; --   +3414700   +5777179
      WHEN 1112 => Ti := "001101001010010011100100010101111101010011010110"; --   +3450084   +5756118
      WHEN 1113 => Ti := "001101010010111010011010010101111000000110111000"; --   +3485338   +5734840
      WHEN 1114 => Ti := "001101011011011111001101010101110010110111000011"; --   +3520461   +5713347
      WHEN 1115 => Ti := "001101100100000001111011010101101101100011110110"; --   +3555451   +5691638
      WHEN 1116 => Ti := "001101101100100010100011010101101000001101010011"; --   +3590307   +5669715
      WHEN 1117 => Ti := "001101110101000001000100010101100010110011011011"; --   +3625028   +5647579
      WHEN 1118 => Ti := "001101111101011101011101010101011101010110001110"; --   +3659613   +5625230
      WHEN 1119 => Ti := "001110000101110111101100010101010111110101101101"; --   +3694060   +5602669
      WHEN 1120 => Ti := "001110001110001111110000010101010010010001111001"; --   +3728368   +5579897
      WHEN 1121 => Ti := "001110010110100101100111010101001100101010110011"; --   +3762535   +5556915
      WHEN 1122 => Ti := "001110011110111001010001010101000111000000011100"; --   +3796561   +5533724
      WHEN 1123 => Ti := "001110100111001010101100010101000001010010110101"; --   +3830444   +5510325
      WHEN 1124 => Ti := "001110101111011001110110010100111011100001111110"; --   +3864182   +5486718
      WHEN 1125 => Ti := "001110110111100110110000010100110101101101111000"; --   +3897776   +5462904
      WHEN 1126 => Ti := "001110111111110001010110010100101111110110100101"; --   +3931222   +5438885
      WHEN 1127 => Ti := "001111000111111001101000010100101001111100000101"; --   +3964520   +5414661
      WHEN 1128 => Ti := "001111001111111111100101010100100011111110011001"; --   +3997669   +5390233
      WHEN 1129 => Ti := "001111011000000011001100010100011101111101100011"; --   +4030668   +5365603
      WHEN 1130 => Ti := "001111100000000100011011010100010111111001100010"; --   +4063515   +5340770
      WHEN 1131 => Ti := "001111101000000011010001010100010001110010011000"; --   +4096209   +5315736
      WHEN 1132 => Ti := "001111101111111111101100010100001011101000000110"; --   +4128748   +5290502
      WHEN 1133 => Ti := "001111110111111001101101010100000101011010101101"; --   +4161133   +5265069
      WHEN 1134 => Ti := "001111111111110001010000010011111111001010001110"; --   +4193360   +5239438
      WHEN 1135 => Ti := "010000000111100110010110010011111000110110101001"; --   +4225430   +5213609
      WHEN 1136 => Ti := "010000001111011000111100010011110010100000000000"; --   +4257340   +5187584
      WHEN 1137 => Ti := "010000010111001001000011010011101100000110010100"; --   +4289091   +5161364
      WHEN 1138 => Ti := "010000011110110110100111010011100101101001100101"; --   +4320679   +5134949
      WHEN 1139 => Ti := "010000100110100001101001010011011111001001110110"; --   +4352105   +5108342
      WHEN 1140 => Ti := "010000101110001010001000010011011000100111000101"; --   +4383368   +5081541
      WHEN 1141 => Ti := "010000110101110000000001010011010010000001010110"; --   +4414465   +5054550
      WHEN 1142 => Ti := "010000111101010011010100010011001011011000101000"; --   +4445396   +5027368
      WHEN 1143 => Ti := "010001000100110100000000010011000100101100111101"; --   +4476160   +4999997
      WHEN 1144 => Ti := "010001001100010010000011010010111101111110010110"; --   +4506755   +4972438
      WHEN 1145 => Ti := "010001010011101101011100010010110111001100110011"; --   +4537180   +4944691
      WHEN 1146 => Ti := "010001011011000110001011010010110000011000010111"; --   +4567435   +4916759
      WHEN 1147 => Ti := "010001100010011100001110010010101001100001000001"; --   +4597518   +4888641
      WHEN 1148 => Ti := "010001101001101111100011010010100010100110110011"; --   +4627427   +4860339
      WHEN 1149 => Ti := "010001110001000000001011010010011011101001101110"; --   +4657163   +4831854
      WHEN 1150 => Ti := "010001111000001110000011010010010100101001110011"; --   +4686723   +4803187
      WHEN 1151 => Ti := "010001111111011001001010010010001101100111000100"; --   +4716106   +4774340
      WHEN 1152 => Ti := "010010000110100001100000010010000110100001100000"; --   +4745312   +4745312
      WHEN 1153 => Ti := "010010001101100111000100010001111111011001001010"; --   +4774340   +4716106
      WHEN 1154 => Ti := "010010010100101001110011010001111000001110000011"; --   +4803187   +4686723
      WHEN 1155 => Ti := "010010011011101001101110010001110001000000001011"; --   +4831854   +4657163
      WHEN 1156 => Ti := "010010100010100110110011010001101001101111100011"; --   +4860339   +4627427
      WHEN 1157 => Ti := "010010101001100001000001010001100010011100001110"; --   +4888641   +4597518
      WHEN 1158 => Ti := "010010110000011000010111010001011011000110001011"; --   +4916759   +4567435
      WHEN 1159 => Ti := "010010110111001100110011010001010011101101011100"; --   +4944691   +4537180
      WHEN 1160 => Ti := "010010111101111110010110010001001100010010000011"; --   +4972438   +4506755
      WHEN 1161 => Ti := "010011000100101100111101010001000100110100000000"; --   +4999997   +4476160
      WHEN 1162 => Ti := "010011001011011000101000010000111101010011010100"; --   +5027368   +4445396
      WHEN 1163 => Ti := "010011010010000001010110010000110101110000000001"; --   +5054550   +4414465
      WHEN 1164 => Ti := "010011011000100111000101010000101110001010001000"; --   +5081541   +4383368
      WHEN 1165 => Ti := "010011011111001001110110010000100110100001101001"; --   +5108342   +4352105
      WHEN 1166 => Ti := "010011100101101001100101010000011110110110100111"; --   +5134949   +4320679
      WHEN 1167 => Ti := "010011101100000110010100010000010111001001000011"; --   +5161364   +4289091
      WHEN 1168 => Ti := "010011110010100000000000010000001111011000111100"; --   +5187584   +4257340
      WHEN 1169 => Ti := "010011111000110110101001010000000111100110010110"; --   +5213609   +4225430
      WHEN 1170 => Ti := "010011111111001010001110001111111111110001010000"; --   +5239438   +4193360
      WHEN 1171 => Ti := "010100000101011010101101001111110111111001101101"; --   +5265069   +4161133
      WHEN 1172 => Ti := "010100001011101000000110001111101111111111101100"; --   +5290502   +4128748
      WHEN 1173 => Ti := "010100010001110010011000001111101000000011010001"; --   +5315736   +4096209
      WHEN 1174 => Ti := "010100010111111001100010001111100000000100011011"; --   +5340770   +4063515
      WHEN 1175 => Ti := "010100011101111101100011001111011000000011001100"; --   +5365603   +4030668
      WHEN 1176 => Ti := "010100100011111110011001001111001111111111100101"; --   +5390233   +3997669
      WHEN 1177 => Ti := "010100101001111100000101001111000111111001101000"; --   +5414661   +3964520
      WHEN 1178 => Ti := "010100101111110110100101001110111111110001010110"; --   +5438885   +3931222
      WHEN 1179 => Ti := "010100110101101101111000001110110111100110110000"; --   +5462904   +3897776
      WHEN 1180 => Ti := "010100111011100001111110001110101111011001110110"; --   +5486718   +3864182
      WHEN 1181 => Ti := "010101000001010010110101001110100111001010101100"; --   +5510325   +3830444
      WHEN 1182 => Ti := "010101000111000000011100001110011110111001010001"; --   +5533724   +3796561
      WHEN 1183 => Ti := "010101001100101010110011001110010110100101100111"; --   +5556915   +3762535
      WHEN 1184 => Ti := "010101010010010001111001001110001110001111110000"; --   +5579897   +3728368
      WHEN 1185 => Ti := "010101010111110101101101001110000101110111101100"; --   +5602669   +3694060
      WHEN 1186 => Ti := "010101011101010110001110001101111101011101011101"; --   +5625230   +3659613
      WHEN 1187 => Ti := "010101100010110011011011001101110101000001000100"; --   +5647579   +3625028
      WHEN 1188 => Ti := "010101101000001101010011001101101100100010100011"; --   +5669715   +3590307
      WHEN 1189 => Ti := "010101101101100011110110001101100100000001111011"; --   +5691638   +3555451
      WHEN 1190 => Ti := "010101110010110111000011001101011011011111001101"; --   +5713347   +3520461
      WHEN 1191 => Ti := "010101111000000110111000001101010010111010011010"; --   +5734840   +3485338
      WHEN 1192 => Ti := "010101111101010011010110001101001010010011100100"; --   +5756118   +3450084
      WHEN 1193 => Ti := "010110000010011100011011001101000001101010101100"; --   +5777179   +3414700
      WHEN 1194 => Ti := "010110000111100010000110001100111000111111110100"; --   +5798022   +3379188
      WHEN 1195 => Ti := "010110001100100100011000001100110000010010111100"; --   +5818648   +3343548
      WHEN 1196 => Ti := "010110010001100011001110001100100111100100000111"; --   +5839054   +3307783
      WHEN 1197 => Ti := "010110010110011110101000001100011110110011010101"; --   +5859240   +3271893
      WHEN 1198 => Ti := "010110011011010110100110001100010110000000101000"; --   +5879206   +3235880
      WHEN 1199 => Ti := "010110100000001011000110001100001101001100000001"; --   +5898950   +3199745
      WHEN 1200 => Ti := "010110100100111100001000001100000100010101100001"; --   +5918472   +3163489
      WHEN 1201 => Ti := "010110101001101001101100001011111011011101001010"; --   +5937772   +3127114
      WHEN 1202 => Ti := "010110101110010011101111001011110010100010111110"; --   +5956847   +3090622
      WHEN 1203 => Ti := "010110110010111010010011001011101001100110111101"; --   +5975699   +3054013
      WHEN 1204 => Ti := "010110110111011101010110001011100000101001001010"; --   +5994326   +3017290
      WHEN 1205 => Ti := "010110111011111100110111001011010111101001100100"; --   +6012727   +2980452
      WHEN 1206 => Ti := "010111000000011000110101001011001110101000001111"; --   +6030901   +2943503
      WHEN 1207 => Ti := "010111000100110001010000001011000101100101001011"; --   +6048848   +2906443
      WHEN 1208 => Ti := "010111001001000110001000001010111100100000011001"; --   +6066568   +2869273
      WHEN 1209 => Ti := "010111001101010111011100001010110011011001111011"; --   +6084060   +2831995
      WHEN 1210 => Ti := "010111010001100101001010001010101010010001110011"; --   +6101322   +2794611
      WHEN 1211 => Ti := "010111010101101111010010001010100001001000000001"; --   +6118354   +2757121
      WHEN 1212 => Ti := "010111011001110101110101001010010111111100101000"; --   +6135157   +2719528
      WHEN 1213 => Ti := "010111011101111000110000001010001110101111101000"; --   +6151728   +2681832
      WHEN 1214 => Ti := "010111100001111000000011001010000101100001000011"; --   +6168067   +2644035
      WHEN 1215 => Ti := "010111100101110011101111001001111100010000111011"; --   +6184175   +2606139
      WHEN 1216 => Ti := "010111101001101011110001001001110010111111010000"; --   +6200049   +2568144
      WHEN 1217 => Ti := "010111101101100000001010001001101001101100000101"; --   +6215690   +2530053
      WHEN 1218 => Ti := "010111110001010000111010001001100000010111011011"; --   +6231098   +2491867
      WHEN 1219 => Ti := "010111110100111101111110001001010111000001010011"; --   +6246270   +2453587
      WHEN 1220 => Ti := "010111111000100111010111001001001101101001101110"; --   +6261207   +2415214
      WHEN 1221 => Ti := "010111111100001101000101001001000100010000101110"; --   +6275909   +2376750
      WHEN 1222 => Ti := "010111111111101111000110001000111010110110010101"; --   +6290374   +2338197
      WHEN 1223 => Ti := "011000000011001101011011001000110001011010100100"; --   +6304603   +2299556
      WHEN 1224 => Ti := "011000000110101000000010001000100111111101011101"; --   +6318594   +2260829
      WHEN 1225 => Ti := "011000001001111110111011001000011110011111000000"; --   +6332347   +2222016
      WHEN 1226 => Ti := "011000001101010010000110001000010100111111010000"; --   +6345862   +2183120
      WHEN 1227 => Ti := "011000010000100001100010001000001011011110001101"; --   +6359138   +2144141
      WHEN 1228 => Ti := "011000010011101101001110001000000001111011111010"; --   +6372174   +2105082
      WHEN 1229 => Ti := "011000010110110101001011000111111000011000010111"; --   +6384971   +2065943
      WHEN 1230 => Ti := "011000011001111001010111000111101110110011100111"; --   +6397527   +2026727
      WHEN 1231 => Ti := "011000011100111001110011000111100101001101101010"; --   +6409843   +1987434
      WHEN 1232 => Ti := "011000011111110110011101000111011011100110100011"; --   +6421917   +1948067
      WHEN 1233 => Ti := "011000100010101111010101000111010001111110010010"; --   +6433749   +1908626
      WHEN 1234 => Ti := "011000100101100100011011000111001000010100111001"; --   +6445339   +1869113
      WHEN 1235 => Ti := "011000101000010101101110000110111110101010011010"; --   +6456686   +1829530
      WHEN 1236 => Ti := "011000101011000011001110000110110100111110110110"; --   +6467790   +1789878
      WHEN 1237 => Ti := "011000101101101100111011000110101011010010001111"; --   +6478651   +1750159
      WHEN 1238 => Ti := "011000110000010010110100000110100001100100100110"; --   +6489268   +1710374
      WHEN 1239 => Ti := "011000110010110100111000000110010111110101111100"; --   +6499640   +1670524
      WHEN 1240 => Ti := "011000110101010011001000000110001110000110010100"; --   +6509768   +1630612
      WHEN 1241 => Ti := "011000110111101101100011000110000100010101101110"; --   +6519651   +1590638
      WHEN 1242 => Ti := "011000111010000100001000000101111010100100001100"; --   +6529288   +1550604
      WHEN 1243 => Ti := "011000111100010110111000000101110000110001110000"; --   +6538680   +1510512
      WHEN 1244 => Ti := "011000111110100101110001000101100110111110011011"; --   +6547825   +1470363
      WHEN 1245 => Ti := "011001000000110000110100000101011101001010001110"; --   +6556724   +1430158
      WHEN 1246 => Ti := "011001000010110111111111000101010011010101001100"; --   +6565375   +1389900
      WHEN 1247 => Ti := "011001000100111011010100000101001001011111010110"; --   +6573780   +1349590
      WHEN 1248 => Ti := "011001000110111010110001000100111111101000101100"; --   +6581937   +1309228
      WHEN 1249 => Ti := "011001001000110110010111000100110101110001010010"; --   +6589847   +1268818
      WHEN 1250 => Ti := "011001001010101110000100000100101011111001000111"; --   +6597508   +1228359
      WHEN 1251 => Ti := "011001001100100001111001000100100010000000001111"; --   +6604921   +1187855
      WHEN 1252 => Ti := "011001001110010001110101000100011000000110101001"; --   +6612085   +1147305
      WHEN 1253 => Ti := "011001001111111101111000000100001110001100011001"; --   +6619000   +1106713
      WHEN 1254 => Ti := "011001010001100110000010000100000100010001011110"; --   +6625666   +1066078
      WHEN 1255 => Ti := "011001010011001010010011000011111010010101111100"; --   +6632083   +1025404
      WHEN 1256 => Ti := "011001010100101010101010000011110000011001110011"; --   +6638250    +984691
      WHEN 1257 => Ti := "011001010110000111000111000011100110011101000101"; --   +6644167    +943941
      WHEN 1258 => Ti := "011001010111011111101010000011011100011111110011"; --   +6649834    +903155
      WHEN 1259 => Ti := "011001011000110100010010000011010010100010000000"; --   +6655250    +862336
      WHEN 1260 => Ti := "011001011010000101000000000011001000100011101100"; --   +6660416    +821484
      WHEN 1261 => Ti := "011001011011010001110011000010111110100100111001"; --   +6665331    +780601
      WHEN 1262 => Ti := "011001011100011010101011000010110100100101101000"; --   +6669995    +739688
      WHEN 1263 => Ti := "011001011101011111101001000010101010100101111100"; --   +6674409    +698748
      WHEN 1264 => Ti := "011001011110100000101010000010100000100101110101"; --   +6678570    +657781
      WHEN 1265 => Ti := "011001011111011101110001000010010110100101010110"; --   +6682481    +616790
      WHEN 1266 => Ti := "011001100000010110111011000010001100100100011111"; --   +6686139    +575775
      WHEN 1267 => Ti := "011001100001001100001010000010000010100011010011"; --   +6689546    +534739
      WHEN 1268 => Ti := "011001100001111101011110000001111000100001110011"; --   +6692702    +493683
      WHEN 1269 => Ti := "011001100010101010110101000001101110100000000000"; --   +6695605    +452608
      WHEN 1270 => Ti := "011001100011010100010000000001100100011101111100"; --   +6698256    +411516
      WHEN 1271 => Ti := "011001100011111001101111000001011010011011101000"; --   +6700655    +370408
      WHEN 1272 => Ti := "011001100100011011010010000001010000011001000111"; --   +6702802    +329287
      WHEN 1273 => Ti := "011001100100111000111000000001000110010110011001"; --   +6704696    +288153
      WHEN 1274 => Ti := "011001100101010010100010000000111100010011100001"; --   +6706338    +247009
      WHEN 1275 => Ti := "011001100101101000001111000000110010010000011111"; --   +6707727    +205855
      WHEN 1276 => Ti := "011001100101111010000000000000101000001101010101"; --   +6708864    +164693
      WHEN 1277 => Ti := "011001100110000111110100000000011110001010000101"; --   +6709748    +123525
      WHEN 1278 => Ti := "011001100110010001101100000000010100000110110000"; --   +6710380     +82352
      WHEN 1279 => Ti := "011001100110010111100111000000001010000011011001"; --   +6710759     +41177
      WHEN 1280 => Ti := "011001100110011001100101000000000000000000000000"; --   +6710885         +0
      WHEN 1281 => Ti := "011001100110010111100111111111110101111100100111"; --   +6710759     -41177
      WHEN 1282 => Ti := "011001100110010001101100111111101011111001010000"; --   +6710380     -82352
      WHEN 1283 => Ti := "011001100110000111110100111111100001110101111011"; --   +6709748    -123525
      WHEN 1284 => Ti := "011001100101111010000000111111010111110010101011"; --   +6708864    -164693
      WHEN 1285 => Ti := "011001100101101000001111111111001101101111100001"; --   +6707727    -205855
      WHEN 1286 => Ti := "011001100101010010100010111111000011101100011111"; --   +6706338    -247009
      WHEN 1287 => Ti := "011001100100111000111000111110111001101001100111"; --   +6704696    -288153
      WHEN 1288 => Ti := "011001100100011011010010111110101111100110111001"; --   +6702802    -329287
      WHEN 1289 => Ti := "011001100011111001101111111110100101100100011000"; --   +6700655    -370408
      WHEN 1290 => Ti := "011001100011010100010000111110011011100010000100"; --   +6698256    -411516
      WHEN 1291 => Ti := "011001100010101010110101111110010001100000000000"; --   +6695605    -452608
      WHEN 1292 => Ti := "011001100001111101011110111110000111011110001101"; --   +6692702    -493683
      WHEN 1293 => Ti := "011001100001001100001010111101111101011100101101"; --   +6689546    -534739
      WHEN 1294 => Ti := "011001100000010110111011111101110011011011100001"; --   +6686139    -575775
      WHEN 1295 => Ti := "011001011111011101110001111101101001011010101010"; --   +6682481    -616790
      WHEN 1296 => Ti := "011001011110100000101010111101011111011010001011"; --   +6678570    -657781
      WHEN 1297 => Ti := "011001011101011111101001111101010101011010000100"; --   +6674409    -698748
      WHEN 1298 => Ti := "011001011100011010101011111101001011011010011000"; --   +6669995    -739688
      WHEN 1299 => Ti := "011001011011010001110011111101000001011011000111"; --   +6665331    -780601
      WHEN 1300 => Ti := "011001011010000101000000111100110111011100010100"; --   +6660416    -821484
      WHEN 1301 => Ti := "011001011000110100010010111100101101011110000000"; --   +6655250    -862336
      WHEN 1302 => Ti := "011001010111011111101010111100100011100000001101"; --   +6649834    -903155
      WHEN 1303 => Ti := "011001010110000111000111111100011001100010111011"; --   +6644167    -943941
      WHEN 1304 => Ti := "011001010100101010101010111100001111100110001101"; --   +6638250    -984691
      WHEN 1305 => Ti := "011001010011001010010011111100000101101010000100"; --   +6632083   -1025404
      WHEN 1306 => Ti := "011001010001100110000010111011111011101110100010"; --   +6625666   -1066078
      WHEN 1307 => Ti := "011001001111111101111000111011110001110011100111"; --   +6619000   -1106713
      WHEN 1308 => Ti := "011001001110010001110101111011100111111001010111"; --   +6612085   -1147305
      WHEN 1309 => Ti := "011001001100100001111001111011011101111111110001"; --   +6604921   -1187855
      WHEN 1310 => Ti := "011001001010101110000100111011010100000110111001"; --   +6597508   -1228359
      WHEN 1311 => Ti := "011001001000110110010111111011001010001110101110"; --   +6589847   -1268818
      WHEN 1312 => Ti := "011001000110111010110001111011000000010111010100"; --   +6581937   -1309228
      WHEN 1313 => Ti := "011001000100111011010100111010110110100000101010"; --   +6573780   -1349590
      WHEN 1314 => Ti := "011001000010110111111111111010101100101010110100"; --   +6565375   -1389900
      WHEN 1315 => Ti := "011001000000110000110100111010100010110101110010"; --   +6556724   -1430158
      WHEN 1316 => Ti := "011000111110100101110001111010011001000001100101"; --   +6547825   -1470363
      WHEN 1317 => Ti := "011000111100010110111000111010001111001110010000"; --   +6538680   -1510512
      WHEN 1318 => Ti := "011000111010000100001000111010000101011011110100"; --   +6529288   -1550604
      WHEN 1319 => Ti := "011000110111101101100011111001111011101010010010"; --   +6519651   -1590638
      WHEN 1320 => Ti := "011000110101010011001000111001110001111001101100"; --   +6509768   -1630612
      WHEN 1321 => Ti := "011000110010110100111000111001101000001010000100"; --   +6499640   -1670524
      WHEN 1322 => Ti := "011000110000010010110100111001011110011011011010"; --   +6489268   -1710374
      WHEN 1323 => Ti := "011000101101101100111011111001010100101101110001"; --   +6478651   -1750159
      WHEN 1324 => Ti := "011000101011000011001110111001001011000001001010"; --   +6467790   -1789878
      WHEN 1325 => Ti := "011000101000010101101110111001000001010101100110"; --   +6456686   -1829530
      WHEN 1326 => Ti := "011000100101100100011011111000110111101011000111"; --   +6445339   -1869113
      WHEN 1327 => Ti := "011000100010101111010101111000101110000001101110"; --   +6433749   -1908626
      WHEN 1328 => Ti := "011000011111110110011101111000100100011001011101"; --   +6421917   -1948067
      WHEN 1329 => Ti := "011000011100111001110011111000011010110010010110"; --   +6409843   -1987434
      WHEN 1330 => Ti := "011000011001111001010111111000010001001100011001"; --   +6397527   -2026727
      WHEN 1331 => Ti := "011000010110110101001011111000000111100111101001"; --   +6384971   -2065943
      WHEN 1332 => Ti := "011000010011101101001110110111111110000100000110"; --   +6372174   -2105082
      WHEN 1333 => Ti := "011000010000100001100010110111110100100001110011"; --   +6359138   -2144141
      WHEN 1334 => Ti := "011000001101010010000110110111101011000000110000"; --   +6345862   -2183120
      WHEN 1335 => Ti := "011000001001111110111011110111100001100001000000"; --   +6332347   -2222016
      WHEN 1336 => Ti := "011000000110101000000010110111011000000010100011"; --   +6318594   -2260829
      WHEN 1337 => Ti := "011000000011001101011011110111001110100101011100"; --   +6304603   -2299556
      WHEN 1338 => Ti := "010111111111101111000110110111000101001001101011"; --   +6290374   -2338197
      WHEN 1339 => Ti := "010111111100001101000101110110111011101111010010"; --   +6275909   -2376750
      WHEN 1340 => Ti := "010111111000100111010111110110110010010110010010"; --   +6261207   -2415214
      WHEN 1341 => Ti := "010111110100111101111110110110101000111110101101"; --   +6246270   -2453587
      WHEN 1342 => Ti := "010111110001010000111010110110011111101000100101"; --   +6231098   -2491867
      WHEN 1343 => Ti := "010111101101100000001010110110010110010011111011"; --   +6215690   -2530053
      WHEN 1344 => Ti := "010111101001101011110001110110001101000000110000"; --   +6200049   -2568144
      WHEN 1345 => Ti := "010111100101110011101111110110000011101111000101"; --   +6184175   -2606139
      WHEN 1346 => Ti := "010111100001111000000011110101111010011110111101"; --   +6168067   -2644035
      WHEN 1347 => Ti := "010111011101111000110000110101110001010000011000"; --   +6151728   -2681832
      WHEN 1348 => Ti := "010111011001110101110101110101101000000011011000"; --   +6135157   -2719528
      WHEN 1349 => Ti := "010111010101101111010010110101011110110111111111"; --   +6118354   -2757121
      WHEN 1350 => Ti := "010111010001100101001010110101010101101110001101"; --   +6101322   -2794611
      WHEN 1351 => Ti := "010111001101010111011100110101001100100110000101"; --   +6084060   -2831995
      WHEN 1352 => Ti := "010111001001000110001000110101000011011111100111"; --   +6066568   -2869273
      WHEN 1353 => Ti := "010111000100110001010000110100111010011010110101"; --   +6048848   -2906443
      WHEN 1354 => Ti := "010111000000011000110101110100110001010111110001"; --   +6030901   -2943503
      WHEN 1355 => Ti := "010110111011111100110111110100101000010110011100"; --   +6012727   -2980452
      WHEN 1356 => Ti := "010110110111011101010110110100011111010110110110"; --   +5994326   -3017290
      WHEN 1357 => Ti := "010110110010111010010011110100010110011001000011"; --   +5975699   -3054013
      WHEN 1358 => Ti := "010110101110010011101111110100001101011101000010"; --   +5956847   -3090622
      WHEN 1359 => Ti := "010110101001101001101100110100000100100010110110"; --   +5937772   -3127114
      WHEN 1360 => Ti := "010110100100111100001000110011111011101010011111"; --   +5918472   -3163489
      WHEN 1361 => Ti := "010110100000001011000110110011110010110011111111"; --   +5898950   -3199745
      WHEN 1362 => Ti := "010110011011010110100110110011101001111111011000"; --   +5879206   -3235880
      WHEN 1363 => Ti := "010110010110011110101000110011100001001100101011"; --   +5859240   -3271893
      WHEN 1364 => Ti := "010110010001100011001110110011011000011011111001"; --   +5839054   -3307783
      WHEN 1365 => Ti := "010110001100100100011000110011001111101101000100"; --   +5818648   -3343548
      WHEN 1366 => Ti := "010110000111100010000110110011000111000000001100"; --   +5798022   -3379188
      WHEN 1367 => Ti := "010110000010011100011011110010111110010101010100"; --   +5777179   -3414700
      WHEN 1368 => Ti := "010101111101010011010110110010110101101100011100"; --   +5756118   -3450084
      WHEN 1369 => Ti := "010101111000000110111000110010101101000101100110"; --   +5734840   -3485338
      WHEN 1370 => Ti := "010101110010110111000011110010100100100000110011"; --   +5713347   -3520461
      WHEN 1371 => Ti := "010101101101100011110110110010011011111110000101"; --   +5691638   -3555451
      WHEN 1372 => Ti := "010101101000001101010011110010010011011101011101"; --   +5669715   -3590307
      WHEN 1373 => Ti := "010101100010110011011011110010001010111110111100"; --   +5647579   -3625028
      WHEN 1374 => Ti := "010101011101010110001110110010000010100010100011"; --   +5625230   -3659613
      WHEN 1375 => Ti := "010101010111110101101101110001111010001000010100"; --   +5602669   -3694060
      WHEN 1376 => Ti := "010101010010010001111001110001110001110000010000"; --   +5579897   -3728368
      WHEN 1377 => Ti := "010101001100101010110011110001101001011010011001"; --   +5556915   -3762535
      WHEN 1378 => Ti := "010101000111000000011100110001100001000110101111"; --   +5533724   -3796561
      WHEN 1379 => Ti := "010101000001010010110101110001011000110101010100"; --   +5510325   -3830444
      WHEN 1380 => Ti := "010100111011100001111110110001010000100110001010"; --   +5486718   -3864182
      WHEN 1381 => Ti := "010100110101101101111000110001001000011001010000"; --   +5462904   -3897776
      WHEN 1382 => Ti := "010100101111110110100101110001000000001110101010"; --   +5438885   -3931222
      WHEN 1383 => Ti := "010100101001111100000101110000111000000110011000"; --   +5414661   -3964520
      WHEN 1384 => Ti := "010100100011111110011001110000110000000000011011"; --   +5390233   -3997669
      WHEN 1385 => Ti := "010100011101111101100011110000100111111100110100"; --   +5365603   -4030668
      WHEN 1386 => Ti := "010100010111111001100010110000011111111011100101"; --   +5340770   -4063515
      WHEN 1387 => Ti := "010100010001110010011000110000010111111100101111"; --   +5315736   -4096209
      WHEN 1388 => Ti := "010100001011101000000110110000010000000000010100"; --   +5290502   -4128748
      WHEN 1389 => Ti := "010100000101011010101101110000001000000110010011"; --   +5265069   -4161133
      WHEN 1390 => Ti := "010011111111001010001110110000000000001110110000"; --   +5239438   -4193360
      WHEN 1391 => Ti := "010011111000110110101001101111111000011001101010"; --   +5213609   -4225430
      WHEN 1392 => Ti := "010011110010100000000000101111110000100111000100"; --   +5187584   -4257340
      WHEN 1393 => Ti := "010011101100000110010100101111101000110110111101"; --   +5161364   -4289091
      WHEN 1394 => Ti := "010011100101101001100101101111100001001001011001"; --   +5134949   -4320679
      WHEN 1395 => Ti := "010011011111001001110110101111011001011110010111"; --   +5108342   -4352105
      WHEN 1396 => Ti := "010011011000100111000101101111010001110101111000"; --   +5081541   -4383368
      WHEN 1397 => Ti := "010011010010000001010110101111001010001111111111"; --   +5054550   -4414465
      WHEN 1398 => Ti := "010011001011011000101000101111000010101100101100"; --   +5027368   -4445396
      WHEN 1399 => Ti := "010011000100101100111101101110111011001100000000"; --   +4999997   -4476160
      WHEN 1400 => Ti := "010010111101111110010110101110110011101101111101"; --   +4972438   -4506755
      WHEN 1401 => Ti := "010010110111001100110011101110101100010010100100"; --   +4944691   -4537180
      WHEN 1402 => Ti := "010010110000011000010111101110100100111001110101"; --   +4916759   -4567435
      WHEN 1403 => Ti := "010010101001100001000001101110011101100011110010"; --   +4888641   -4597518
      WHEN 1404 => Ti := "010010100010100110110011101110010110010000011101"; --   +4860339   -4627427
      WHEN 1405 => Ti := "010010011011101001101110101110001110111111110101"; --   +4831854   -4657163
      WHEN 1406 => Ti := "010010010100101001110011101110000111110001111101"; --   +4803187   -4686723
      WHEN 1407 => Ti := "010010001101100111000100101110000000100110110110"; --   +4774340   -4716106
      WHEN 1408 => Ti := "010010000110100001100000101101111001011110100000"; --   +4745312   -4745312
      WHEN 1409 => Ti := "010001111111011001001010101101110010011000111100"; --   +4716106   -4774340
      WHEN 1410 => Ti := "010001111000001110000011101101101011010110001101"; --   +4686723   -4803187
      WHEN 1411 => Ti := "010001110001000000001011101101100100010110010010"; --   +4657163   -4831854
      WHEN 1412 => Ti := "010001101001101111100011101101011101011001001101"; --   +4627427   -4860339
      WHEN 1413 => Ti := "010001100010011100001110101101010110011110111111"; --   +4597518   -4888641
      WHEN 1414 => Ti := "010001011011000110001011101101001111100111101001"; --   +4567435   -4916759
      WHEN 1415 => Ti := "010001010011101101011100101101001000110011001101"; --   +4537180   -4944691
      WHEN 1416 => Ti := "010001001100010010000011101101000010000001101010"; --   +4506755   -4972438
      WHEN 1417 => Ti := "010001000100110100000000101100111011010011000011"; --   +4476160   -4999997
      WHEN 1418 => Ti := "010000111101010011010100101100110100100111011000"; --   +4445396   -5027368
      WHEN 1419 => Ti := "010000110101110000000001101100101101111110101010"; --   +4414465   -5054550
      WHEN 1420 => Ti := "010000101110001010001000101100100111011000111011"; --   +4383368   -5081541
      WHEN 1421 => Ti := "010000100110100001101001101100100000110110001010"; --   +4352105   -5108342
      WHEN 1422 => Ti := "010000011110110110100111101100011010010110011011"; --   +4320679   -5134949
      WHEN 1423 => Ti := "010000010111001001000011101100010011111001101100"; --   +4289091   -5161364
      WHEN 1424 => Ti := "010000001111011000111100101100001101100000000000"; --   +4257340   -5187584
      WHEN 1425 => Ti := "010000000111100110010110101100000111001001010111"; --   +4225430   -5213609
      WHEN 1426 => Ti := "001111111111110001010000101100000000110101110010"; --   +4193360   -5239438
      WHEN 1427 => Ti := "001111110111111001101101101011111010100101010011"; --   +4161133   -5265069
      WHEN 1428 => Ti := "001111101111111111101100101011110100010111111010"; --   +4128748   -5290502
      WHEN 1429 => Ti := "001111101000000011010001101011101110001101101000"; --   +4096209   -5315736
      WHEN 1430 => Ti := "001111100000000100011011101011101000000110011110"; --   +4063515   -5340770
      WHEN 1431 => Ti := "001111011000000011001100101011100010000010011101"; --   +4030668   -5365603
      WHEN 1432 => Ti := "001111001111111111100101101011011100000001100111"; --   +3997669   -5390233
      WHEN 1433 => Ti := "001111000111111001101000101011010110000011111011"; --   +3964520   -5414661
      WHEN 1434 => Ti := "001110111111110001010110101011010000001001011011"; --   +3931222   -5438885
      WHEN 1435 => Ti := "001110110111100110110000101011001010010010001000"; --   +3897776   -5462904
      WHEN 1436 => Ti := "001110101111011001110110101011000100011110000010"; --   +3864182   -5486718
      WHEN 1437 => Ti := "001110100111001010101100101010111110101101001011"; --   +3830444   -5510325
      WHEN 1438 => Ti := "001110011110111001010001101010111000111111100100"; --   +3796561   -5533724
      WHEN 1439 => Ti := "001110010110100101100111101010110011010101001101"; --   +3762535   -5556915
      WHEN 1440 => Ti := "001110001110001111110000101010101101101110000111"; --   +3728368   -5579897
      WHEN 1441 => Ti := "001110000101110111101100101010101000001010010011"; --   +3694060   -5602669
      WHEN 1442 => Ti := "001101111101011101011101101010100010101001110010"; --   +3659613   -5625230
      WHEN 1443 => Ti := "001101110101000001000100101010011101001100100101"; --   +3625028   -5647579
      WHEN 1444 => Ti := "001101101100100010100011101010010111110010101101"; --   +3590307   -5669715
      WHEN 1445 => Ti := "001101100100000001111011101010010010011100001010"; --   +3555451   -5691638
      WHEN 1446 => Ti := "001101011011011111001101101010001101001000111101"; --   +3520461   -5713347
      WHEN 1447 => Ti := "001101010010111010011010101010000111111001001000"; --   +3485338   -5734840
      WHEN 1448 => Ti := "001101001010010011100100101010000010101100101010"; --   +3450084   -5756118
      WHEN 1449 => Ti := "001101000001101010101100101001111101100011100101"; --   +3414700   -5777179
      WHEN 1450 => Ti := "001100111000111111110100101001111000011101111010"; --   +3379188   -5798022
      WHEN 1451 => Ti := "001100110000010010111100101001110011011011101000"; --   +3343548   -5818648
      WHEN 1452 => Ti := "001100100111100100000111101001101110011100110010"; --   +3307783   -5839054
      WHEN 1453 => Ti := "001100011110110011010101101001101001100001011000"; --   +3271893   -5859240
      WHEN 1454 => Ti := "001100010110000000101000101001100100101001011010"; --   +3235880   -5879206
      WHEN 1455 => Ti := "001100001101001100000001101001011111110100111010"; --   +3199745   -5898950
      WHEN 1456 => Ti := "001100000100010101100001101001011011000011111000"; --   +3163489   -5918472
      WHEN 1457 => Ti := "001011111011011101001010101001010110010110010100"; --   +3127114   -5937772
      WHEN 1458 => Ti := "001011110010100010111110101001010001101100010001"; --   +3090622   -5956847
      WHEN 1459 => Ti := "001011101001100110111101101001001101000101101101"; --   +3054013   -5975699
      WHEN 1460 => Ti := "001011100000101001001010101001001000100010101010"; --   +3017290   -5994326
      WHEN 1461 => Ti := "001011010111101001100100101001000100000011001001"; --   +2980452   -6012727
      WHEN 1462 => Ti := "001011001110101000001111101000111111100111001011"; --   +2943503   -6030901
      WHEN 1463 => Ti := "001011000101100101001011101000111011001110110000"; --   +2906443   -6048848
      WHEN 1464 => Ti := "001010111100100000011001101000110110111001111000"; --   +2869273   -6066568
      WHEN 1465 => Ti := "001010110011011001111011101000110010101000100100"; --   +2831995   -6084060
      WHEN 1466 => Ti := "001010101010010001110011101000101110011010110110"; --   +2794611   -6101322
      WHEN 1467 => Ti := "001010100001001000000001101000101010010000101110"; --   +2757121   -6118354
      WHEN 1468 => Ti := "001010010111111100101000101000100110001010001011"; --   +2719528   -6135157
      WHEN 1469 => Ti := "001010001110101111101000101000100010000111010000"; --   +2681832   -6151728
      WHEN 1470 => Ti := "001010000101100001000011101000011110000111111101"; --   +2644035   -6168067
      WHEN 1471 => Ti := "001001111100010000111011101000011010001100010001"; --   +2606139   -6184175
      WHEN 1472 => Ti := "001001110010111111010000101000010110010100001111"; --   +2568144   -6200049
      WHEN 1473 => Ti := "001001101001101100000101101000010010011111110110"; --   +2530053   -6215690
      WHEN 1474 => Ti := "001001100000010111011011101000001110101111000110"; --   +2491867   -6231098
      WHEN 1475 => Ti := "001001010111000001010011101000001011000010000010"; --   +2453587   -6246270
      WHEN 1476 => Ti := "001001001101101001101110101000000111011000101001"; --   +2415214   -6261207
      WHEN 1477 => Ti := "001001000100010000101110101000000011110010111011"; --   +2376750   -6275909
      WHEN 1478 => Ti := "001000111010110110010101101000000000010000111010"; --   +2338197   -6290374
      WHEN 1479 => Ti := "001000110001011010100100100111111100110010100101"; --   +2299556   -6304603
      WHEN 1480 => Ti := "001000100111111101011101100111111001010111111110"; --   +2260829   -6318594
      WHEN 1481 => Ti := "001000011110011111000000100111110110000001000101"; --   +2222016   -6332347
      WHEN 1482 => Ti := "001000010100111111010000100111110010101101111010"; --   +2183120   -6345862
      WHEN 1483 => Ti := "001000001011011110001101100111101111011110011110"; --   +2144141   -6359138
      WHEN 1484 => Ti := "001000000001111011111010100111101100010010110010"; --   +2105082   -6372174
      WHEN 1485 => Ti := "000111111000011000010111100111101001001010110101"; --   +2065943   -6384971
      WHEN 1486 => Ti := "000111101110110011100111100111100110000110101001"; --   +2026727   -6397527
      WHEN 1487 => Ti := "000111100101001101101010100111100011000110001101"; --   +1987434   -6409843
      WHEN 1488 => Ti := "000111011011100110100011100111100000001001100011"; --   +1948067   -6421917
      WHEN 1489 => Ti := "000111010001111110010010100111011101010000101011"; --   +1908626   -6433749
      WHEN 1490 => Ti := "000111001000010100111001100111011010011011100101"; --   +1869113   -6445339
      WHEN 1491 => Ti := "000110111110101010011010100111010111101010010010"; --   +1829530   -6456686
      WHEN 1492 => Ti := "000110110100111110110110100111010100111100110010"; --   +1789878   -6467790
      WHEN 1493 => Ti := "000110101011010010001111100111010010010011000101"; --   +1750159   -6478651
      WHEN 1494 => Ti := "000110100001100100100110100111001111101101001100"; --   +1710374   -6489268
      WHEN 1495 => Ti := "000110010111110101111100100111001101001011001000"; --   +1670524   -6499640
      WHEN 1496 => Ti := "000110001110000110010100100111001010101100111000"; --   +1630612   -6509768
      WHEN 1497 => Ti := "000110000100010101101110100111001000010010011101"; --   +1590638   -6519651
      WHEN 1498 => Ti := "000101111010100100001100100111000101111011111000"; --   +1550604   -6529288
      WHEN 1499 => Ti := "000101110000110001110000100111000011101001001000"; --   +1510512   -6538680
      WHEN 1500 => Ti := "000101100110111110011011100111000001011010001111"; --   +1470363   -6547825
      WHEN 1501 => Ti := "000101011101001010001110100110111111001111001100"; --   +1430158   -6556724
      WHEN 1502 => Ti := "000101010011010101001100100110111101001000000001"; --   +1389900   -6565375
      WHEN 1503 => Ti := "000101001001011111010110100110111011000100101100"; --   +1349590   -6573780
      WHEN 1504 => Ti := "000100111111101000101100100110111001000101001111"; --   +1309228   -6581937
      WHEN 1505 => Ti := "000100110101110001010010100110110111001001101001"; --   +1268818   -6589847
      WHEN 1506 => Ti := "000100101011111001000111100110110101010001111100"; --   +1228359   -6597508
      WHEN 1507 => Ti := "000100100010000000001111100110110011011110000111"; --   +1187855   -6604921
      WHEN 1508 => Ti := "000100011000000110101001100110110001101110001011"; --   +1147305   -6612085
      WHEN 1509 => Ti := "000100001110001100011001100110110000000010001000"; --   +1106713   -6619000
      WHEN 1510 => Ti := "000100000100010001011110100110101110011001111110"; --   +1066078   -6625666
      WHEN 1511 => Ti := "000011111010010101111100100110101100110101101101"; --   +1025404   -6632083
      WHEN 1512 => Ti := "000011110000011001110011100110101011010101010110"; --    +984691   -6638250
      WHEN 1513 => Ti := "000011100110011101000101100110101001111000111001"; --    +943941   -6644167
      WHEN 1514 => Ti := "000011011100011111110011100110101000100000010110"; --    +903155   -6649834
      WHEN 1515 => Ti := "000011010010100010000000100110100111001011101110"; --    +862336   -6655250
      WHEN 1516 => Ti := "000011001000100011101100100110100101111011000000"; --    +821484   -6660416
      WHEN 1517 => Ti := "000010111110100100111001100110100100101110001101"; --    +780601   -6665331
      WHEN 1518 => Ti := "000010110100100101101000100110100011100101010101"; --    +739688   -6669995
      WHEN 1519 => Ti := "000010101010100101111100100110100010100000010111"; --    +698748   -6674409
      WHEN 1520 => Ti := "000010100000100101110101100110100001011111010110"; --    +657781   -6678570
      WHEN 1521 => Ti := "000010010110100101010110100110100000100010001111"; --    +616790   -6682481
      WHEN 1522 => Ti := "000010001100100100011111100110011111101001000101"; --    +575775   -6686139
      WHEN 1523 => Ti := "000010000010100011010011100110011110110011110110"; --    +534739   -6689546
      WHEN 1524 => Ti := "000001111000100001110011100110011110000010100010"; --    +493683   -6692702
      WHEN 1525 => Ti := "000001101110100000000000100110011101010101001011"; --    +452608   -6695605
      WHEN 1526 => Ti := "000001100100011101111100100110011100101011110000"; --    +411516   -6698256
      WHEN 1527 => Ti := "000001011010011011101000100110011100000110010001"; --    +370408   -6700655
      WHEN 1528 => Ti := "000001010000011001000111100110011011100100101110"; --    +329287   -6702802
      WHEN 1529 => Ti := "000001000110010110011001100110011011000111001000"; --    +288153   -6704696
      WHEN 1530 => Ti := "000000111100010011100001100110011010101101011110"; --    +247009   -6706338
      WHEN 1531 => Ti := "000000110010010000011111100110011010010111110001"; --    +205855   -6707727
      WHEN 1532 => Ti := "000000101000001101010101100110011010000110000000"; --    +164693   -6708864
      WHEN 1533 => Ti := "000000011110001010000101100110011001111000001100"; --    +123525   -6709748
      WHEN 1534 => Ti := "000000010100000110110000100110011001101110010100"; --     +82352   -6710380
      WHEN 1535 => Ti := "000000001010000011011001100110011001101000011001"; --     +41177   -6710759
      WHEN 1536 => Ti := "000000000000000000000000100110011001100110011011"; --         +0   -6710885
      WHEN 1537 => Ti := "111111110101111100100111100110011001101000011001"; --     -41177   -6710759
      WHEN 1538 => Ti := "111111101011111001010000100110011001101110010100"; --     -82352   -6710380
      WHEN 1539 => Ti := "111111100001110101111011100110011001111000001100"; --    -123525   -6709748
      WHEN 1540 => Ti := "111111010111110010101011100110011010000110000000"; --    -164693   -6708864
      WHEN 1541 => Ti := "111111001101101111100001100110011010010111110001"; --    -205855   -6707727
      WHEN 1542 => Ti := "111111000011101100011111100110011010101101011110"; --    -247009   -6706338
      WHEN 1543 => Ti := "111110111001101001100111100110011011000111001000"; --    -288153   -6704696
      WHEN 1544 => Ti := "111110101111100110111001100110011011100100101110"; --    -329287   -6702802
      WHEN 1545 => Ti := "111110100101100100011000100110011100000110010001"; --    -370408   -6700655
      WHEN 1546 => Ti := "111110011011100010000100100110011100101011110000"; --    -411516   -6698256
      WHEN 1547 => Ti := "111110010001100000000000100110011101010101001011"; --    -452608   -6695605
      WHEN 1548 => Ti := "111110000111011110001101100110011110000010100010"; --    -493683   -6692702
      WHEN 1549 => Ti := "111101111101011100101101100110011110110011110110"; --    -534739   -6689546
      WHEN 1550 => Ti := "111101110011011011100001100110011111101001000101"; --    -575775   -6686139
      WHEN 1551 => Ti := "111101101001011010101010100110100000100010001111"; --    -616790   -6682481
      WHEN 1552 => Ti := "111101011111011010001011100110100001011111010110"; --    -657781   -6678570
      WHEN 1553 => Ti := "111101010101011010000100100110100010100000010111"; --    -698748   -6674409
      WHEN 1554 => Ti := "111101001011011010011000100110100011100101010101"; --    -739688   -6669995
      WHEN 1555 => Ti := "111101000001011011000111100110100100101110001101"; --    -780601   -6665331
      WHEN 1556 => Ti := "111100110111011100010100100110100101111011000000"; --    -821484   -6660416
      WHEN 1557 => Ti := "111100101101011110000000100110100111001011101110"; --    -862336   -6655250
      WHEN 1558 => Ti := "111100100011100000001101100110101000100000010110"; --    -903155   -6649834
      WHEN 1559 => Ti := "111100011001100010111011100110101001111000111001"; --    -943941   -6644167
      WHEN 1560 => Ti := "111100001111100110001101100110101011010101010110"; --    -984691   -6638250
      WHEN 1561 => Ti := "111100000101101010000100100110101100110101101101"; --   -1025404   -6632083
      WHEN 1562 => Ti := "111011111011101110100010100110101110011001111110"; --   -1066078   -6625666
      WHEN 1563 => Ti := "111011110001110011100111100110110000000010001000"; --   -1106713   -6619000
      WHEN 1564 => Ti := "111011100111111001010111100110110001101110001011"; --   -1147305   -6612085
      WHEN 1565 => Ti := "111011011101111111110001100110110011011110000111"; --   -1187855   -6604921
      WHEN 1566 => Ti := "111011010100000110111001100110110101010001111100"; --   -1228359   -6597508
      WHEN 1567 => Ti := "111011001010001110101110100110110111001001101001"; --   -1268818   -6589847
      WHEN 1568 => Ti := "111011000000010111010100100110111001000101001111"; --   -1309228   -6581937
      WHEN 1569 => Ti := "111010110110100000101010100110111011000100101100"; --   -1349590   -6573780
      WHEN 1570 => Ti := "111010101100101010110100100110111101001000000001"; --   -1389900   -6565375
      WHEN 1571 => Ti := "111010100010110101110010100110111111001111001100"; --   -1430158   -6556724
      WHEN 1572 => Ti := "111010011001000001100101100111000001011010001111"; --   -1470363   -6547825
      WHEN 1573 => Ti := "111010001111001110010000100111000011101001001000"; --   -1510512   -6538680
      WHEN 1574 => Ti := "111010000101011011110100100111000101111011111000"; --   -1550604   -6529288
      WHEN 1575 => Ti := "111001111011101010010010100111001000010010011101"; --   -1590638   -6519651
      WHEN 1576 => Ti := "111001110001111001101100100111001010101100111000"; --   -1630612   -6509768
      WHEN 1577 => Ti := "111001101000001010000100100111001101001011001000"; --   -1670524   -6499640
      WHEN 1578 => Ti := "111001011110011011011010100111001111101101001100"; --   -1710374   -6489268
      WHEN 1579 => Ti := "111001010100101101110001100111010010010011000101"; --   -1750159   -6478651
      WHEN 1580 => Ti := "111001001011000001001010100111010100111100110010"; --   -1789878   -6467790
      WHEN 1581 => Ti := "111001000001010101100110100111010111101010010010"; --   -1829530   -6456686
      WHEN 1582 => Ti := "111000110111101011000111100111011010011011100101"; --   -1869113   -6445339
      WHEN 1583 => Ti := "111000101110000001101110100111011101010000101011"; --   -1908626   -6433749
      WHEN 1584 => Ti := "111000100100011001011101100111100000001001100011"; --   -1948067   -6421917
      WHEN 1585 => Ti := "111000011010110010010110100111100011000110001101"; --   -1987434   -6409843
      WHEN 1586 => Ti := "111000010001001100011001100111100110000110101001"; --   -2026727   -6397527
      WHEN 1587 => Ti := "111000000111100111101001100111101001001010110101"; --   -2065943   -6384971
      WHEN 1588 => Ti := "110111111110000100000110100111101100010010110010"; --   -2105082   -6372174
      WHEN 1589 => Ti := "110111110100100001110011100111101111011110011110"; --   -2144141   -6359138
      WHEN 1590 => Ti := "110111101011000000110000100111110010101101111010"; --   -2183120   -6345862
      WHEN 1591 => Ti := "110111100001100001000000100111110110000001000101"; --   -2222016   -6332347
      WHEN 1592 => Ti := "110111011000000010100011100111111001010111111110"; --   -2260829   -6318594
      WHEN 1593 => Ti := "110111001110100101011100100111111100110010100101"; --   -2299556   -6304603
      WHEN 1594 => Ti := "110111000101001001101011101000000000010000111010"; --   -2338197   -6290374
      WHEN 1595 => Ti := "110110111011101111010010101000000011110010111011"; --   -2376750   -6275909
      WHEN 1596 => Ti := "110110110010010110010010101000000111011000101001"; --   -2415214   -6261207
      WHEN 1597 => Ti := "110110101000111110101101101000001011000010000010"; --   -2453587   -6246270
      WHEN 1598 => Ti := "110110011111101000100101101000001110101111000110"; --   -2491867   -6231098
      WHEN 1599 => Ti := "110110010110010011111011101000010010011111110110"; --   -2530053   -6215690
      WHEN 1600 => Ti := "110110001101000000110000101000010110010100001111"; --   -2568144   -6200049
      WHEN 1601 => Ti := "110110000011101111000101101000011010001100010001"; --   -2606139   -6184175
      WHEN 1602 => Ti := "110101111010011110111101101000011110000111111101"; --   -2644035   -6168067
      WHEN 1603 => Ti := "110101110001010000011000101000100010000111010000"; --   -2681832   -6151728
      WHEN 1604 => Ti := "110101101000000011011000101000100110001010001011"; --   -2719528   -6135157
      WHEN 1605 => Ti := "110101011110110111111111101000101010010000101110"; --   -2757121   -6118354
      WHEN 1606 => Ti := "110101010101101110001101101000101110011010110110"; --   -2794611   -6101322
      WHEN 1607 => Ti := "110101001100100110000101101000110010101000100100"; --   -2831995   -6084060
      WHEN 1608 => Ti := "110101000011011111100111101000110110111001111000"; --   -2869273   -6066568
      WHEN 1609 => Ti := "110100111010011010110101101000111011001110110000"; --   -2906443   -6048848
      WHEN 1610 => Ti := "110100110001010111110001101000111111100111001011"; --   -2943503   -6030901
      WHEN 1611 => Ti := "110100101000010110011100101001000100000011001001"; --   -2980452   -6012727
      WHEN 1612 => Ti := "110100011111010110110110101001001000100010101010"; --   -3017290   -5994326
      WHEN 1613 => Ti := "110100010110011001000011101001001101000101101101"; --   -3054013   -5975699
      WHEN 1614 => Ti := "110100001101011101000010101001010001101100010001"; --   -3090622   -5956847
      WHEN 1615 => Ti := "110100000100100010110110101001010110010110010100"; --   -3127114   -5937772
      WHEN 1616 => Ti := "110011111011101010011111101001011011000011111000"; --   -3163489   -5918472
      WHEN 1617 => Ti := "110011110010110011111111101001011111110100111010"; --   -3199745   -5898950
      WHEN 1618 => Ti := "110011101001111111011000101001100100101001011010"; --   -3235880   -5879206
      WHEN 1619 => Ti := "110011100001001100101011101001101001100001011000"; --   -3271893   -5859240
      WHEN 1620 => Ti := "110011011000011011111001101001101110011100110010"; --   -3307783   -5839054
      WHEN 1621 => Ti := "110011001111101101000100101001110011011011101000"; --   -3343548   -5818648
      WHEN 1622 => Ti := "110011000111000000001100101001111000011101111010"; --   -3379188   -5798022
      WHEN 1623 => Ti := "110010111110010101010100101001111101100011100101"; --   -3414700   -5777179
      WHEN 1624 => Ti := "110010110101101100011100101010000010101100101010"; --   -3450084   -5756118
      WHEN 1625 => Ti := "110010101101000101100110101010000111111001001000"; --   -3485338   -5734840
      WHEN 1626 => Ti := "110010100100100000110011101010001101001000111101"; --   -3520461   -5713347
      WHEN 1627 => Ti := "110010011011111110000101101010010010011100001010"; --   -3555451   -5691638
      WHEN 1628 => Ti := "110010010011011101011101101010010111110010101101"; --   -3590307   -5669715
      WHEN 1629 => Ti := "110010001010111110111100101010011101001100100101"; --   -3625028   -5647579
      WHEN 1630 => Ti := "110010000010100010100011101010100010101001110010"; --   -3659613   -5625230
      WHEN 1631 => Ti := "110001111010001000010100101010101000001010010011"; --   -3694060   -5602669
      WHEN 1632 => Ti := "110001110001110000010000101010101101101110000111"; --   -3728368   -5579897
      WHEN 1633 => Ti := "110001101001011010011001101010110011010101001101"; --   -3762535   -5556915
      WHEN 1634 => Ti := "110001100001000110101111101010111000111111100100"; --   -3796561   -5533724
      WHEN 1635 => Ti := "110001011000110101010100101010111110101101001011"; --   -3830444   -5510325
      WHEN 1636 => Ti := "110001010000100110001010101011000100011110000010"; --   -3864182   -5486718
      WHEN 1637 => Ti := "110001001000011001010000101011001010010010001000"; --   -3897776   -5462904
      WHEN 1638 => Ti := "110001000000001110101010101011010000001001011011"; --   -3931222   -5438885
      WHEN 1639 => Ti := "110000111000000110011000101011010110000011111011"; --   -3964520   -5414661
      WHEN 1640 => Ti := "110000110000000000011011101011011100000001100111"; --   -3997669   -5390233
      WHEN 1641 => Ti := "110000100111111100110100101011100010000010011101"; --   -4030668   -5365603
      WHEN 1642 => Ti := "110000011111111011100101101011101000000110011110"; --   -4063515   -5340770
      WHEN 1643 => Ti := "110000010111111100101111101011101110001101101000"; --   -4096209   -5315736
      WHEN 1644 => Ti := "110000010000000000010100101011110100010111111010"; --   -4128748   -5290502
      WHEN 1645 => Ti := "110000001000000110010011101011111010100101010011"; --   -4161133   -5265069
      WHEN 1646 => Ti := "110000000000001110110000101100000000110101110010"; --   -4193360   -5239438
      WHEN 1647 => Ti := "101111111000011001101010101100000111001001010111"; --   -4225430   -5213609
      WHEN 1648 => Ti := "101111110000100111000100101100001101100000000000"; --   -4257340   -5187584
      WHEN 1649 => Ti := "101111101000110110111101101100010011111001101100"; --   -4289091   -5161364
      WHEN 1650 => Ti := "101111100001001001011001101100011010010110011011"; --   -4320679   -5134949
      WHEN 1651 => Ti := "101111011001011110010111101100100000110110001010"; --   -4352105   -5108342
      WHEN 1652 => Ti := "101111010001110101111000101100100111011000111011"; --   -4383368   -5081541
      WHEN 1653 => Ti := "101111001010001111111111101100101101111110101010"; --   -4414465   -5054550
      WHEN 1654 => Ti := "101111000010101100101100101100110100100111011000"; --   -4445396   -5027368
      WHEN 1655 => Ti := "101110111011001100000000101100111011010011000011"; --   -4476160   -4999997
      WHEN 1656 => Ti := "101110110011101101111101101101000010000001101010"; --   -4506755   -4972438
      WHEN 1657 => Ti := "101110101100010010100100101101001000110011001101"; --   -4537180   -4944691
      WHEN 1658 => Ti := "101110100100111001110101101101001111100111101001"; --   -4567435   -4916759
      WHEN 1659 => Ti := "101110011101100011110010101101010110011110111111"; --   -4597518   -4888641
      WHEN 1660 => Ti := "101110010110010000011101101101011101011001001101"; --   -4627427   -4860339
      WHEN 1661 => Ti := "101110001110111111110101101101100100010110010010"; --   -4657163   -4831854
      WHEN 1662 => Ti := "101110000111110001111101101101101011010110001101"; --   -4686723   -4803187
      WHEN 1663 => Ti := "101110000000100110110110101101110010011000111100"; --   -4716106   -4774340
      WHEN 1664 => Ti := "101101111001011110100000101101111001011110100000"; --   -4745312   -4745312
      WHEN 1665 => Ti := "101101110010011000111100101110000000100110110110"; --   -4774340   -4716106
      WHEN 1666 => Ti := "101101101011010110001101101110000111110001111101"; --   -4803187   -4686723
      WHEN 1667 => Ti := "101101100100010110010010101110001110111111110101"; --   -4831854   -4657163
      WHEN 1668 => Ti := "101101011101011001001101101110010110010000011101"; --   -4860339   -4627427
      WHEN 1669 => Ti := "101101010110011110111111101110011101100011110010"; --   -4888641   -4597518
      WHEN 1670 => Ti := "101101001111100111101001101110100100111001110101"; --   -4916759   -4567435
      WHEN 1671 => Ti := "101101001000110011001101101110101100010010100100"; --   -4944691   -4537180
      WHEN 1672 => Ti := "101101000010000001101010101110110011101101111101"; --   -4972438   -4506755
      WHEN 1673 => Ti := "101100111011010011000011101110111011001100000000"; --   -4999997   -4476160
      WHEN 1674 => Ti := "101100110100100111011000101111000010101100101100"; --   -5027368   -4445396
      WHEN 1675 => Ti := "101100101101111110101010101111001010001111111111"; --   -5054550   -4414465
      WHEN 1676 => Ti := "101100100111011000111011101111010001110101111000"; --   -5081541   -4383368
      WHEN 1677 => Ti := "101100100000110110001010101111011001011110010111"; --   -5108342   -4352105
      WHEN 1678 => Ti := "101100011010010110011011101111100001001001011001"; --   -5134949   -4320679
      WHEN 1679 => Ti := "101100010011111001101100101111101000110110111101"; --   -5161364   -4289091
      WHEN 1680 => Ti := "101100001101100000000000101111110000100111000100"; --   -5187584   -4257340
      WHEN 1681 => Ti := "101100000111001001010111101111111000011001101010"; --   -5213609   -4225430
      WHEN 1682 => Ti := "101100000000110101110010110000000000001110110000"; --   -5239438   -4193360
      WHEN 1683 => Ti := "101011111010100101010011110000001000000110010011"; --   -5265069   -4161133
      WHEN 1684 => Ti := "101011110100010111111010110000010000000000010100"; --   -5290502   -4128748
      WHEN 1685 => Ti := "101011101110001101101000110000010111111100101111"; --   -5315736   -4096209
      WHEN 1686 => Ti := "101011101000000110011110110000011111111011100101"; --   -5340770   -4063515
      WHEN 1687 => Ti := "101011100010000010011101110000100111111100110100"; --   -5365603   -4030668
      WHEN 1688 => Ti := "101011011100000001100111110000110000000000011011"; --   -5390233   -3997669
      WHEN 1689 => Ti := "101011010110000011111011110000111000000110011000"; --   -5414661   -3964520
      WHEN 1690 => Ti := "101011010000001001011011110001000000001110101010"; --   -5438885   -3931222
      WHEN 1691 => Ti := "101011001010010010001000110001001000011001010000"; --   -5462904   -3897776
      WHEN 1692 => Ti := "101011000100011110000010110001010000100110001010"; --   -5486718   -3864182
      WHEN 1693 => Ti := "101010111110101101001011110001011000110101010100"; --   -5510325   -3830444
      WHEN 1694 => Ti := "101010111000111111100100110001100001000110101111"; --   -5533724   -3796561
      WHEN 1695 => Ti := "101010110011010101001101110001101001011010011001"; --   -5556915   -3762535
      WHEN 1696 => Ti := "101010101101101110000111110001110001110000010000"; --   -5579897   -3728368
      WHEN 1697 => Ti := "101010101000001010010011110001111010001000010100"; --   -5602669   -3694060
      WHEN 1698 => Ti := "101010100010101001110010110010000010100010100011"; --   -5625230   -3659613
      WHEN 1699 => Ti := "101010011101001100100101110010001010111110111100"; --   -5647579   -3625028
      WHEN 1700 => Ti := "101010010111110010101101110010010011011101011101"; --   -5669715   -3590307
      WHEN 1701 => Ti := "101010010010011100001010110010011011111110000101"; --   -5691638   -3555451
      WHEN 1702 => Ti := "101010001101001000111101110010100100100000110011"; --   -5713347   -3520461
      WHEN 1703 => Ti := "101010000111111001001000110010101101000101100110"; --   -5734840   -3485338
      WHEN 1704 => Ti := "101010000010101100101010110010110101101100011100"; --   -5756118   -3450084
      WHEN 1705 => Ti := "101001111101100011100101110010111110010101010100"; --   -5777179   -3414700
      WHEN 1706 => Ti := "101001111000011101111010110011000111000000001100"; --   -5798022   -3379188
      WHEN 1707 => Ti := "101001110011011011101000110011001111101101000100"; --   -5818648   -3343548
      WHEN 1708 => Ti := "101001101110011100110010110011011000011011111001"; --   -5839054   -3307783
      WHEN 1709 => Ti := "101001101001100001011000110011100001001100101011"; --   -5859240   -3271893
      WHEN 1710 => Ti := "101001100100101001011010110011101001111111011000"; --   -5879206   -3235880
      WHEN 1711 => Ti := "101001011111110100111010110011110010110011111111"; --   -5898950   -3199745
      WHEN 1712 => Ti := "101001011011000011111000110011111011101010011111"; --   -5918472   -3163489
      WHEN 1713 => Ti := "101001010110010110010100110100000100100010110110"; --   -5937772   -3127114
      WHEN 1714 => Ti := "101001010001101100010001110100001101011101000010"; --   -5956847   -3090622
      WHEN 1715 => Ti := "101001001101000101101101110100010110011001000011"; --   -5975699   -3054013
      WHEN 1716 => Ti := "101001001000100010101010110100011111010110110110"; --   -5994326   -3017290
      WHEN 1717 => Ti := "101001000100000011001001110100101000010110011100"; --   -6012727   -2980452
      WHEN 1718 => Ti := "101000111111100111001011110100110001010111110001"; --   -6030901   -2943503
      WHEN 1719 => Ti := "101000111011001110110000110100111010011010110101"; --   -6048848   -2906443
      WHEN 1720 => Ti := "101000110110111001111000110101000011011111100111"; --   -6066568   -2869273
      WHEN 1721 => Ti := "101000110010101000100100110101001100100110000101"; --   -6084060   -2831995
      WHEN 1722 => Ti := "101000101110011010110110110101010101101110001101"; --   -6101322   -2794611
      WHEN 1723 => Ti := "101000101010010000101110110101011110110111111111"; --   -6118354   -2757121
      WHEN 1724 => Ti := "101000100110001010001011110101101000000011011000"; --   -6135157   -2719528
      WHEN 1725 => Ti := "101000100010000111010000110101110001010000011000"; --   -6151728   -2681832
      WHEN 1726 => Ti := "101000011110000111111101110101111010011110111101"; --   -6168067   -2644035
      WHEN 1727 => Ti := "101000011010001100010001110110000011101111000101"; --   -6184175   -2606139
      WHEN 1728 => Ti := "101000010110010100001111110110001101000000110000"; --   -6200049   -2568144
      WHEN 1729 => Ti := "101000010010011111110110110110010110010011111011"; --   -6215690   -2530053
      WHEN 1730 => Ti := "101000001110101111000110110110011111101000100101"; --   -6231098   -2491867
      WHEN 1731 => Ti := "101000001011000010000010110110101000111110101101"; --   -6246270   -2453587
      WHEN 1732 => Ti := "101000000111011000101001110110110010010110010010"; --   -6261207   -2415214
      WHEN 1733 => Ti := "101000000011110010111011110110111011101111010010"; --   -6275909   -2376750
      WHEN 1734 => Ti := "101000000000010000111010110111000101001001101011"; --   -6290374   -2338197
      WHEN 1735 => Ti := "100111111100110010100101110111001110100101011100"; --   -6304603   -2299556
      WHEN 1736 => Ti := "100111111001010111111110110111011000000010100011"; --   -6318594   -2260829
      WHEN 1737 => Ti := "100111110110000001000101110111100001100001000000"; --   -6332347   -2222016
      WHEN 1738 => Ti := "100111110010101101111010110111101011000000110000"; --   -6345862   -2183120
      WHEN 1739 => Ti := "100111101111011110011110110111110100100001110011"; --   -6359138   -2144141
      WHEN 1740 => Ti := "100111101100010010110010110111111110000100000110"; --   -6372174   -2105082
      WHEN 1741 => Ti := "100111101001001010110101111000000111100111101001"; --   -6384971   -2065943
      WHEN 1742 => Ti := "100111100110000110101001111000010001001100011001"; --   -6397527   -2026727
      WHEN 1743 => Ti := "100111100011000110001101111000011010110010010110"; --   -6409843   -1987434
      WHEN 1744 => Ti := "100111100000001001100011111000100100011001011101"; --   -6421917   -1948067
      WHEN 1745 => Ti := "100111011101010000101011111000101110000001101110"; --   -6433749   -1908626
      WHEN 1746 => Ti := "100111011010011011100101111000110111101011000111"; --   -6445339   -1869113
      WHEN 1747 => Ti := "100111010111101010010010111001000001010101100110"; --   -6456686   -1829530
      WHEN 1748 => Ti := "100111010100111100110010111001001011000001001010"; --   -6467790   -1789878
      WHEN 1749 => Ti := "100111010010010011000101111001010100101101110001"; --   -6478651   -1750159
      WHEN 1750 => Ti := "100111001111101101001100111001011110011011011010"; --   -6489268   -1710374
      WHEN 1751 => Ti := "100111001101001011001000111001101000001010000100"; --   -6499640   -1670524
      WHEN 1752 => Ti := "100111001010101100111000111001110001111001101100"; --   -6509768   -1630612
      WHEN 1753 => Ti := "100111001000010010011101111001111011101010010010"; --   -6519651   -1590638
      WHEN 1754 => Ti := "100111000101111011111000111010000101011011110100"; --   -6529288   -1550604
      WHEN 1755 => Ti := "100111000011101001001000111010001111001110010000"; --   -6538680   -1510512
      WHEN 1756 => Ti := "100111000001011010001111111010011001000001100101"; --   -6547825   -1470363
      WHEN 1757 => Ti := "100110111111001111001100111010100010110101110010"; --   -6556724   -1430158
      WHEN 1758 => Ti := "100110111101001000000001111010101100101010110100"; --   -6565375   -1389900
      WHEN 1759 => Ti := "100110111011000100101100111010110110100000101010"; --   -6573780   -1349590
      WHEN 1760 => Ti := "100110111001000101001111111011000000010111010100"; --   -6581937   -1309228
      WHEN 1761 => Ti := "100110110111001001101001111011001010001110101110"; --   -6589847   -1268818
      WHEN 1762 => Ti := "100110110101010001111100111011010100000110111001"; --   -6597508   -1228359
      WHEN 1763 => Ti := "100110110011011110000111111011011101111111110001"; --   -6604921   -1187855
      WHEN 1764 => Ti := "100110110001101110001011111011100111111001010111"; --   -6612085   -1147305
      WHEN 1765 => Ti := "100110110000000010001000111011110001110011100111"; --   -6619000   -1106713
      WHEN 1766 => Ti := "100110101110011001111110111011111011101110100010"; --   -6625666   -1066078
      WHEN 1767 => Ti := "100110101100110101101101111100000101101010000100"; --   -6632083   -1025404
      WHEN 1768 => Ti := "100110101011010101010110111100001111100110001101"; --   -6638250    -984691
      WHEN 1769 => Ti := "100110101001111000111001111100011001100010111011"; --   -6644167    -943941
      WHEN 1770 => Ti := "100110101000100000010110111100100011100000001101"; --   -6649834    -903155
      WHEN 1771 => Ti := "100110100111001011101110111100101101011110000000"; --   -6655250    -862336
      WHEN 1772 => Ti := "100110100101111011000000111100110111011100010100"; --   -6660416    -821484
      WHEN 1773 => Ti := "100110100100101110001101111101000001011011000111"; --   -6665331    -780601
      WHEN 1774 => Ti := "100110100011100101010101111101001011011010011000"; --   -6669995    -739688
      WHEN 1775 => Ti := "100110100010100000010111111101010101011010000100"; --   -6674409    -698748
      WHEN 1776 => Ti := "100110100001011111010110111101011111011010001011"; --   -6678570    -657781
      WHEN 1777 => Ti := "100110100000100010001111111101101001011010101010"; --   -6682481    -616790
      WHEN 1778 => Ti := "100110011111101001000101111101110011011011100001"; --   -6686139    -575775
      WHEN 1779 => Ti := "100110011110110011110110111101111101011100101101"; --   -6689546    -534739
      WHEN 1780 => Ti := "100110011110000010100010111110000111011110001101"; --   -6692702    -493683
      WHEN 1781 => Ti := "100110011101010101001011111110010001100000000000"; --   -6695605    -452608
      WHEN 1782 => Ti := "100110011100101011110000111110011011100010000100"; --   -6698256    -411516
      WHEN 1783 => Ti := "100110011100000110010001111110100101100100011000"; --   -6700655    -370408
      WHEN 1784 => Ti := "100110011011100100101110111110101111100110111001"; --   -6702802    -329287
      WHEN 1785 => Ti := "100110011011000111001000111110111001101001100111"; --   -6704696    -288153
      WHEN 1786 => Ti := "100110011010101101011110111111000011101100011111"; --   -6706338    -247009
      WHEN 1787 => Ti := "100110011010010111110001111111001101101111100001"; --   -6707727    -205855
      WHEN 1788 => Ti := "100110011010000110000000111111010111110010101011"; --   -6708864    -164693
      WHEN 1789 => Ti := "100110011001111000001100111111100001110101111011"; --   -6709748    -123525
      WHEN 1790 => Ti := "100110011001101110010100111111101011111001010000"; --   -6710380     -82352
      WHEN 1791 => Ti := "100110011001101000011001111111110101111100100111"; --   -6710759     -41177
      WHEN 1792 => Ti := "100110011001100110011011000000000000000000000000"; --   -6710885         +0
      WHEN 1793 => Ti := "100110011001101000011001000000001010000011011001"; --   -6710759     +41177
      WHEN 1794 => Ti := "100110011001101110010100000000010100000110110000"; --   -6710380     +82352
      WHEN 1795 => Ti := "100110011001111000001100000000011110001010000101"; --   -6709748    +123525
      WHEN 1796 => Ti := "100110011010000110000000000000101000001101010101"; --   -6708864    +164693
      WHEN 1797 => Ti := "100110011010010111110001000000110010010000011111"; --   -6707727    +205855
      WHEN 1798 => Ti := "100110011010101101011110000000111100010011100001"; --   -6706338    +247009
      WHEN 1799 => Ti := "100110011011000111001000000001000110010110011001"; --   -6704696    +288153
      WHEN 1800 => Ti := "100110011011100100101110000001010000011001000111"; --   -6702802    +329287
      WHEN 1801 => Ti := "100110011100000110010001000001011010011011101000"; --   -6700655    +370408
      WHEN 1802 => Ti := "100110011100101011110000000001100100011101111100"; --   -6698256    +411516
      WHEN 1803 => Ti := "100110011101010101001011000001101110100000000000"; --   -6695605    +452608
      WHEN 1804 => Ti := "100110011110000010100010000001111000100001110011"; --   -6692702    +493683
      WHEN 1805 => Ti := "100110011110110011110110000010000010100011010011"; --   -6689546    +534739
      WHEN 1806 => Ti := "100110011111101001000101000010001100100100011111"; --   -6686139    +575775
      WHEN 1807 => Ti := "100110100000100010001111000010010110100101010110"; --   -6682481    +616790
      WHEN 1808 => Ti := "100110100001011111010110000010100000100101110101"; --   -6678570    +657781
      WHEN 1809 => Ti := "100110100010100000010111000010101010100101111100"; --   -6674409    +698748
      WHEN 1810 => Ti := "100110100011100101010101000010110100100101101000"; --   -6669995    +739688
      WHEN 1811 => Ti := "100110100100101110001101000010111110100100111001"; --   -6665331    +780601
      WHEN 1812 => Ti := "100110100101111011000000000011001000100011101100"; --   -6660416    +821484
      WHEN 1813 => Ti := "100110100111001011101110000011010010100010000000"; --   -6655250    +862336
      WHEN 1814 => Ti := "100110101000100000010110000011011100011111110011"; --   -6649834    +903155
      WHEN 1815 => Ti := "100110101001111000111001000011100110011101000101"; --   -6644167    +943941
      WHEN 1816 => Ti := "100110101011010101010110000011110000011001110011"; --   -6638250    +984691
      WHEN 1817 => Ti := "100110101100110101101101000011111010010101111100"; --   -6632083   +1025404
      WHEN 1818 => Ti := "100110101110011001111110000100000100010001011110"; --   -6625666   +1066078
      WHEN 1819 => Ti := "100110110000000010001000000100001110001100011001"; --   -6619000   +1106713
      WHEN 1820 => Ti := "100110110001101110001011000100011000000110101001"; --   -6612085   +1147305
      WHEN 1821 => Ti := "100110110011011110000111000100100010000000001111"; --   -6604921   +1187855
      WHEN 1822 => Ti := "100110110101010001111100000100101011111001000111"; --   -6597508   +1228359
      WHEN 1823 => Ti := "100110110111001001101001000100110101110001010010"; --   -6589847   +1268818
      WHEN 1824 => Ti := "100110111001000101001111000100111111101000101100"; --   -6581937   +1309228
      WHEN 1825 => Ti := "100110111011000100101100000101001001011111010110"; --   -6573780   +1349590
      WHEN 1826 => Ti := "100110111101001000000001000101010011010101001100"; --   -6565375   +1389900
      WHEN 1827 => Ti := "100110111111001111001100000101011101001010001110"; --   -6556724   +1430158
      WHEN 1828 => Ti := "100111000001011010001111000101100110111110011011"; --   -6547825   +1470363
      WHEN 1829 => Ti := "100111000011101001001000000101110000110001110000"; --   -6538680   +1510512
      WHEN 1830 => Ti := "100111000101111011111000000101111010100100001100"; --   -6529288   +1550604
      WHEN 1831 => Ti := "100111001000010010011101000110000100010101101110"; --   -6519651   +1590638
      WHEN 1832 => Ti := "100111001010101100111000000110001110000110010100"; --   -6509768   +1630612
      WHEN 1833 => Ti := "100111001101001011001000000110010111110101111100"; --   -6499640   +1670524
      WHEN 1834 => Ti := "100111001111101101001100000110100001100100100110"; --   -6489268   +1710374
      WHEN 1835 => Ti := "100111010010010011000101000110101011010010001111"; --   -6478651   +1750159
      WHEN 1836 => Ti := "100111010100111100110010000110110100111110110110"; --   -6467790   +1789878
      WHEN 1837 => Ti := "100111010111101010010010000110111110101010011010"; --   -6456686   +1829530
      WHEN 1838 => Ti := "100111011010011011100101000111001000010100111001"; --   -6445339   +1869113
      WHEN 1839 => Ti := "100111011101010000101011000111010001111110010010"; --   -6433749   +1908626
      WHEN 1840 => Ti := "100111100000001001100011000111011011100110100011"; --   -6421917   +1948067
      WHEN 1841 => Ti := "100111100011000110001101000111100101001101101010"; --   -6409843   +1987434
      WHEN 1842 => Ti := "100111100110000110101001000111101110110011100111"; --   -6397527   +2026727
      WHEN 1843 => Ti := "100111101001001010110101000111111000011000010111"; --   -6384971   +2065943
      WHEN 1844 => Ti := "100111101100010010110010001000000001111011111010"; --   -6372174   +2105082
      WHEN 1845 => Ti := "100111101111011110011110001000001011011110001101"; --   -6359138   +2144141
      WHEN 1846 => Ti := "100111110010101101111010001000010100111111010000"; --   -6345862   +2183120
      WHEN 1847 => Ti := "100111110110000001000101001000011110011111000000"; --   -6332347   +2222016
      WHEN 1848 => Ti := "100111111001010111111110001000100111111101011101"; --   -6318594   +2260829
      WHEN 1849 => Ti := "100111111100110010100101001000110001011010100100"; --   -6304603   +2299556
      WHEN 1850 => Ti := "101000000000010000111010001000111010110110010101"; --   -6290374   +2338197
      WHEN 1851 => Ti := "101000000011110010111011001001000100010000101110"; --   -6275909   +2376750
      WHEN 1852 => Ti := "101000000111011000101001001001001101101001101110"; --   -6261207   +2415214
      WHEN 1853 => Ti := "101000001011000010000010001001010111000001010011"; --   -6246270   +2453587
      WHEN 1854 => Ti := "101000001110101111000110001001100000010111011011"; --   -6231098   +2491867
      WHEN 1855 => Ti := "101000010010011111110110001001101001101100000101"; --   -6215690   +2530053
      WHEN 1856 => Ti := "101000010110010100001111001001110010111111010000"; --   -6200049   +2568144
      WHEN 1857 => Ti := "101000011010001100010001001001111100010000111011"; --   -6184175   +2606139
      WHEN 1858 => Ti := "101000011110000111111101001010000101100001000011"; --   -6168067   +2644035
      WHEN 1859 => Ti := "101000100010000111010000001010001110101111101000"; --   -6151728   +2681832
      WHEN 1860 => Ti := "101000100110001010001011001010010111111100101000"; --   -6135157   +2719528
      WHEN 1861 => Ti := "101000101010010000101110001010100001001000000001"; --   -6118354   +2757121
      WHEN 1862 => Ti := "101000101110011010110110001010101010010001110011"; --   -6101322   +2794611
      WHEN 1863 => Ti := "101000110010101000100100001010110011011001111011"; --   -6084060   +2831995
      WHEN 1864 => Ti := "101000110110111001111000001010111100100000011001"; --   -6066568   +2869273
      WHEN 1865 => Ti := "101000111011001110110000001011000101100101001011"; --   -6048848   +2906443
      WHEN 1866 => Ti := "101000111111100111001011001011001110101000001111"; --   -6030901   +2943503
      WHEN 1867 => Ti := "101001000100000011001001001011010111101001100100"; --   -6012727   +2980452
      WHEN 1868 => Ti := "101001001000100010101010001011100000101001001010"; --   -5994326   +3017290
      WHEN 1869 => Ti := "101001001101000101101101001011101001100110111101"; --   -5975699   +3054013
      WHEN 1870 => Ti := "101001010001101100010001001011110010100010111110"; --   -5956847   +3090622
      WHEN 1871 => Ti := "101001010110010110010100001011111011011101001010"; --   -5937772   +3127114
      WHEN 1872 => Ti := "101001011011000011111000001100000100010101100001"; --   -5918472   +3163489
      WHEN 1873 => Ti := "101001011111110100111010001100001101001100000001"; --   -5898950   +3199745
      WHEN 1874 => Ti := "101001100100101001011010001100010110000000101000"; --   -5879206   +3235880
      WHEN 1875 => Ti := "101001101001100001011000001100011110110011010101"; --   -5859240   +3271893
      WHEN 1876 => Ti := "101001101110011100110010001100100111100100000111"; --   -5839054   +3307783
      WHEN 1877 => Ti := "101001110011011011101000001100110000010010111100"; --   -5818648   +3343548
      WHEN 1878 => Ti := "101001111000011101111010001100111000111111110100"; --   -5798022   +3379188
      WHEN 1879 => Ti := "101001111101100011100101001101000001101010101100"; --   -5777179   +3414700
      WHEN 1880 => Ti := "101010000010101100101010001101001010010011100100"; --   -5756118   +3450084
      WHEN 1881 => Ti := "101010000111111001001000001101010010111010011010"; --   -5734840   +3485338
      WHEN 1882 => Ti := "101010001101001000111101001101011011011111001101"; --   -5713347   +3520461
      WHEN 1883 => Ti := "101010010010011100001010001101100100000001111011"; --   -5691638   +3555451
      WHEN 1884 => Ti := "101010010111110010101101001101101100100010100011"; --   -5669715   +3590307
      WHEN 1885 => Ti := "101010011101001100100101001101110101000001000100"; --   -5647579   +3625028
      WHEN 1886 => Ti := "101010100010101001110010001101111101011101011101"; --   -5625230   +3659613
      WHEN 1887 => Ti := "101010101000001010010011001110000101110111101100"; --   -5602669   +3694060
      WHEN 1888 => Ti := "101010101101101110000111001110001110001111110000"; --   -5579897   +3728368
      WHEN 1889 => Ti := "101010110011010101001101001110010110100101100111"; --   -5556915   +3762535
      WHEN 1890 => Ti := "101010111000111111100100001110011110111001010001"; --   -5533724   +3796561
      WHEN 1891 => Ti := "101010111110101101001011001110100111001010101100"; --   -5510325   +3830444
      WHEN 1892 => Ti := "101011000100011110000010001110101111011001110110"; --   -5486718   +3864182
      WHEN 1893 => Ti := "101011001010010010001000001110110111100110110000"; --   -5462904   +3897776
      WHEN 1894 => Ti := "101011010000001001011011001110111111110001010110"; --   -5438885   +3931222
      WHEN 1895 => Ti := "101011010110000011111011001111000111111001101000"; --   -5414661   +3964520
      WHEN 1896 => Ti := "101011011100000001100111001111001111111111100101"; --   -5390233   +3997669
      WHEN 1897 => Ti := "101011100010000010011101001111011000000011001100"; --   -5365603   +4030668
      WHEN 1898 => Ti := "101011101000000110011110001111100000000100011011"; --   -5340770   +4063515
      WHEN 1899 => Ti := "101011101110001101101000001111101000000011010001"; --   -5315736   +4096209
      WHEN 1900 => Ti := "101011110100010111111010001111101111111111101100"; --   -5290502   +4128748
      WHEN 1901 => Ti := "101011111010100101010011001111110111111001101101"; --   -5265069   +4161133
      WHEN 1902 => Ti := "101100000000110101110010001111111111110001010000"; --   -5239438   +4193360
      WHEN 1903 => Ti := "101100000111001001010111010000000111100110010110"; --   -5213609   +4225430
      WHEN 1904 => Ti := "101100001101100000000000010000001111011000111100"; --   -5187584   +4257340
      WHEN 1905 => Ti := "101100010011111001101100010000010111001001000011"; --   -5161364   +4289091
      WHEN 1906 => Ti := "101100011010010110011011010000011110110110100111"; --   -5134949   +4320679
      WHEN 1907 => Ti := "101100100000110110001010010000100110100001101001"; --   -5108342   +4352105
      WHEN 1908 => Ti := "101100100111011000111011010000101110001010001000"; --   -5081541   +4383368
      WHEN 1909 => Ti := "101100101101111110101010010000110101110000000001"; --   -5054550   +4414465
      WHEN 1910 => Ti := "101100110100100111011000010000111101010011010100"; --   -5027368   +4445396
      WHEN 1911 => Ti := "101100111011010011000011010001000100110100000000"; --   -4999997   +4476160
      WHEN 1912 => Ti := "101101000010000001101010010001001100010010000011"; --   -4972438   +4506755
      WHEN 1913 => Ti := "101101001000110011001101010001010011101101011100"; --   -4944691   +4537180
      WHEN 1914 => Ti := "101101001111100111101001010001011011000110001011"; --   -4916759   +4567435
      WHEN 1915 => Ti := "101101010110011110111111010001100010011100001110"; --   -4888641   +4597518
      WHEN 1916 => Ti := "101101011101011001001101010001101001101111100011"; --   -4860339   +4627427
      WHEN 1917 => Ti := "101101100100010110010010010001110001000000001011"; --   -4831854   +4657163
      WHEN 1918 => Ti := "101101101011010110001101010001111000001110000011"; --   -4803187   +4686723
      WHEN 1919 => Ti := "101101110010011000111100010001111111011001001010"; --   -4774340   +4716106
      WHEN 1920 => Ti := "101101111001011110100000010010000110100001100000"; --   -4745312   +4745312
      WHEN 1921 => Ti := "101110000000100110110110010010001101100111000100"; --   -4716106   +4774340
      WHEN 1922 => Ti := "101110000111110001111101010010010100101001110011"; --   -4686723   +4803187
      WHEN 1923 => Ti := "101110001110111111110101010010011011101001101110"; --   -4657163   +4831854
      WHEN 1924 => Ti := "101110010110010000011101010010100010100110110011"; --   -4627427   +4860339
      WHEN 1925 => Ti := "101110011101100011110010010010101001100001000001"; --   -4597518   +4888641
      WHEN 1926 => Ti := "101110100100111001110101010010110000011000010111"; --   -4567435   +4916759
      WHEN 1927 => Ti := "101110101100010010100100010010110111001100110011"; --   -4537180   +4944691
      WHEN 1928 => Ti := "101110110011101101111101010010111101111110010110"; --   -4506755   +4972438
      WHEN 1929 => Ti := "101110111011001100000000010011000100101100111101"; --   -4476160   +4999997
      WHEN 1930 => Ti := "101111000010101100101100010011001011011000101000"; --   -4445396   +5027368
      WHEN 1931 => Ti := "101111001010001111111111010011010010000001010110"; --   -4414465   +5054550
      WHEN 1932 => Ti := "101111010001110101111000010011011000100111000101"; --   -4383368   +5081541
      WHEN 1933 => Ti := "101111011001011110010111010011011111001001110110"; --   -4352105   +5108342
      WHEN 1934 => Ti := "101111100001001001011001010011100101101001100101"; --   -4320679   +5134949
      WHEN 1935 => Ti := "101111101000110110111101010011101100000110010100"; --   -4289091   +5161364
      WHEN 1936 => Ti := "101111110000100111000100010011110010100000000000"; --   -4257340   +5187584
      WHEN 1937 => Ti := "101111111000011001101010010011111000110110101001"; --   -4225430   +5213609
      WHEN 1938 => Ti := "110000000000001110110000010011111111001010001110"; --   -4193360   +5239438
      WHEN 1939 => Ti := "110000001000000110010011010100000101011010101101"; --   -4161133   +5265069
      WHEN 1940 => Ti := "110000010000000000010100010100001011101000000110"; --   -4128748   +5290502
      WHEN 1941 => Ti := "110000010111111100101111010100010001110010011000"; --   -4096209   +5315736
      WHEN 1942 => Ti := "110000011111111011100101010100010111111001100010"; --   -4063515   +5340770
      WHEN 1943 => Ti := "110000100111111100110100010100011101111101100011"; --   -4030668   +5365603
      WHEN 1944 => Ti := "110000110000000000011011010100100011111110011001"; --   -3997669   +5390233
      WHEN 1945 => Ti := "110000111000000110011000010100101001111100000101"; --   -3964520   +5414661
      WHEN 1946 => Ti := "110001000000001110101010010100101111110110100101"; --   -3931222   +5438885
      WHEN 1947 => Ti := "110001001000011001010000010100110101101101111000"; --   -3897776   +5462904
      WHEN 1948 => Ti := "110001010000100110001010010100111011100001111110"; --   -3864182   +5486718
      WHEN 1949 => Ti := "110001011000110101010100010101000001010010110101"; --   -3830444   +5510325
      WHEN 1950 => Ti := "110001100001000110101111010101000111000000011100"; --   -3796561   +5533724
      WHEN 1951 => Ti := "110001101001011010011001010101001100101010110011"; --   -3762535   +5556915
      WHEN 1952 => Ti := "110001110001110000010000010101010010010001111001"; --   -3728368   +5579897
      WHEN 1953 => Ti := "110001111010001000010100010101010111110101101101"; --   -3694060   +5602669
      WHEN 1954 => Ti := "110010000010100010100011010101011101010110001110"; --   -3659613   +5625230
      WHEN 1955 => Ti := "110010001010111110111100010101100010110011011011"; --   -3625028   +5647579
      WHEN 1956 => Ti := "110010010011011101011101010101101000001101010011"; --   -3590307   +5669715
      WHEN 1957 => Ti := "110010011011111110000101010101101101100011110110"; --   -3555451   +5691638
      WHEN 1958 => Ti := "110010100100100000110011010101110010110111000011"; --   -3520461   +5713347
      WHEN 1959 => Ti := "110010101101000101100110010101111000000110111000"; --   -3485338   +5734840
      WHEN 1960 => Ti := "110010110101101100011100010101111101010011010110"; --   -3450084   +5756118
      WHEN 1961 => Ti := "110010111110010101010100010110000010011100011011"; --   -3414700   +5777179
      WHEN 1962 => Ti := "110011000111000000001100010110000111100010000110"; --   -3379188   +5798022
      WHEN 1963 => Ti := "110011001111101101000100010110001100100100011000"; --   -3343548   +5818648
      WHEN 1964 => Ti := "110011011000011011111001010110010001100011001110"; --   -3307783   +5839054
      WHEN 1965 => Ti := "110011100001001100101011010110010110011110101000"; --   -3271893   +5859240
      WHEN 1966 => Ti := "110011101001111111011000010110011011010110100110"; --   -3235880   +5879206
      WHEN 1967 => Ti := "110011110010110011111111010110100000001011000110"; --   -3199745   +5898950
      WHEN 1968 => Ti := "110011111011101010011111010110100100111100001000"; --   -3163489   +5918472
      WHEN 1969 => Ti := "110100000100100010110110010110101001101001101100"; --   -3127114   +5937772
      WHEN 1970 => Ti := "110100001101011101000010010110101110010011101111"; --   -3090622   +5956847
      WHEN 1971 => Ti := "110100010110011001000011010110110010111010010011"; --   -3054013   +5975699
      WHEN 1972 => Ti := "110100011111010110110110010110110111011101010110"; --   -3017290   +5994326
      WHEN 1973 => Ti := "110100101000010110011100010110111011111100110111"; --   -2980452   +6012727
      WHEN 1974 => Ti := "110100110001010111110001010111000000011000110101"; --   -2943503   +6030901
      WHEN 1975 => Ti := "110100111010011010110101010111000100110001010000"; --   -2906443   +6048848
      WHEN 1976 => Ti := "110101000011011111100111010111001001000110001000"; --   -2869273   +6066568
      WHEN 1977 => Ti := "110101001100100110000101010111001101010111011100"; --   -2831995   +6084060
      WHEN 1978 => Ti := "110101010101101110001101010111010001100101001010"; --   -2794611   +6101322
      WHEN 1979 => Ti := "110101011110110111111111010111010101101111010010"; --   -2757121   +6118354
      WHEN 1980 => Ti := "110101101000000011011000010111011001110101110101"; --   -2719528   +6135157
      WHEN 1981 => Ti := "110101110001010000011000010111011101111000110000"; --   -2681832   +6151728
      WHEN 1982 => Ti := "110101111010011110111101010111100001111000000011"; --   -2644035   +6168067
      WHEN 1983 => Ti := "110110000011101111000101010111100101110011101111"; --   -2606139   +6184175
      WHEN 1984 => Ti := "110110001101000000110000010111101001101011110001"; --   -2568144   +6200049
      WHEN 1985 => Ti := "110110010110010011111011010111101101100000001010"; --   -2530053   +6215690
      WHEN 1986 => Ti := "110110011111101000100101010111110001010000111010"; --   -2491867   +6231098
      WHEN 1987 => Ti := "110110101000111110101101010111110100111101111110"; --   -2453587   +6246270
      WHEN 1988 => Ti := "110110110010010110010010010111111000100111010111"; --   -2415214   +6261207
      WHEN 1989 => Ti := "110110111011101111010010010111111100001101000101"; --   -2376750   +6275909
      WHEN 1990 => Ti := "110111000101001001101011010111111111101111000110"; --   -2338197   +6290374
      WHEN 1991 => Ti := "110111001110100101011100011000000011001101011011"; --   -2299556   +6304603
      WHEN 1992 => Ti := "110111011000000010100011011000000110101000000010"; --   -2260829   +6318594
      WHEN 1993 => Ti := "110111100001100001000000011000001001111110111011"; --   -2222016   +6332347
      WHEN 1994 => Ti := "110111101011000000110000011000001101010010000110"; --   -2183120   +6345862
      WHEN 1995 => Ti := "110111110100100001110011011000010000100001100010"; --   -2144141   +6359138
      WHEN 1996 => Ti := "110111111110000100000110011000010011101101001110"; --   -2105082   +6372174
      WHEN 1997 => Ti := "111000000111100111101001011000010110110101001011"; --   -2065943   +6384971
      WHEN 1998 => Ti := "111000010001001100011001011000011001111001010111"; --   -2026727   +6397527
      WHEN 1999 => Ti := "111000011010110010010110011000011100111001110011"; --   -1987434   +6409843
      WHEN 2000 => Ti := "111000100100011001011101011000011111110110011101"; --   -1948067   +6421917
      WHEN 2001 => Ti := "111000101110000001101110011000100010101111010101"; --   -1908626   +6433749
      WHEN 2002 => Ti := "111000110111101011000111011000100101100100011011"; --   -1869113   +6445339
      WHEN 2003 => Ti := "111001000001010101100110011000101000010101101110"; --   -1829530   +6456686
      WHEN 2004 => Ti := "111001001011000001001010011000101011000011001110"; --   -1789878   +6467790
      WHEN 2005 => Ti := "111001010100101101110001011000101101101100111011"; --   -1750159   +6478651
      WHEN 2006 => Ti := "111001011110011011011010011000110000010010110100"; --   -1710374   +6489268
      WHEN 2007 => Ti := "111001101000001010000100011000110010110100111000"; --   -1670524   +6499640
      WHEN 2008 => Ti := "111001110001111001101100011000110101010011001000"; --   -1630612   +6509768
      WHEN 2009 => Ti := "111001111011101010010010011000110111101101100011"; --   -1590638   +6519651
      WHEN 2010 => Ti := "111010000101011011110100011000111010000100001000"; --   -1550604   +6529288
      WHEN 2011 => Ti := "111010001111001110010000011000111100010110111000"; --   -1510512   +6538680
      WHEN 2012 => Ti := "111010011001000001100101011000111110100101110001"; --   -1470363   +6547825
      WHEN 2013 => Ti := "111010100010110101110010011001000000110000110100"; --   -1430158   +6556724
      WHEN 2014 => Ti := "111010101100101010110100011001000010110111111111"; --   -1389900   +6565375
      WHEN 2015 => Ti := "111010110110100000101010011001000100111011010100"; --   -1349590   +6573780
      WHEN 2016 => Ti := "111011000000010111010100011001000110111010110001"; --   -1309228   +6581937
      WHEN 2017 => Ti := "111011001010001110101110011001001000110110010111"; --   -1268818   +6589847
      WHEN 2018 => Ti := "111011010100000110111001011001001010101110000100"; --   -1228359   +6597508
      WHEN 2019 => Ti := "111011011101111111110001011001001100100001111001"; --   -1187855   +6604921
      WHEN 2020 => Ti := "111011100111111001010111011001001110010001110101"; --   -1147305   +6612085
      WHEN 2021 => Ti := "111011110001110011100111011001001111111101111000"; --   -1106713   +6619000
      WHEN 2022 => Ti := "111011111011101110100010011001010001100110000010"; --   -1066078   +6625666
      WHEN 2023 => Ti := "111100000101101010000100011001010011001010010011"; --   -1025404   +6632083
      WHEN 2024 => Ti := "111100001111100110001101011001010100101010101010"; --    -984691   +6638250
      WHEN 2025 => Ti := "111100011001100010111011011001010110000111000111"; --    -943941   +6644167
      WHEN 2026 => Ti := "111100100011100000001101011001010111011111101010"; --    -903155   +6649834
      WHEN 2027 => Ti := "111100101101011110000000011001011000110100010010"; --    -862336   +6655250
      WHEN 2028 => Ti := "111100110111011100010100011001011010000101000000"; --    -821484   +6660416
      WHEN 2029 => Ti := "111101000001011011000111011001011011010001110011"; --    -780601   +6665331
      WHEN 2030 => Ti := "111101001011011010011000011001011100011010101011"; --    -739688   +6669995
      WHEN 2031 => Ti := "111101010101011010000100011001011101011111101001"; --    -698748   +6674409
      WHEN 2032 => Ti := "111101011111011010001011011001011110100000101010"; --    -657781   +6678570
      WHEN 2033 => Ti := "111101101001011010101010011001011111011101110001"; --    -616790   +6682481
      WHEN 2034 => Ti := "111101110011011011100001011001100000010110111011"; --    -575775   +6686139
      WHEN 2035 => Ti := "111101111101011100101101011001100001001100001010"; --    -534739   +6689546
      WHEN 2036 => Ti := "111110000111011110001101011001100001111101011110"; --    -493683   +6692702
      WHEN 2037 => Ti := "111110010001100000000000011001100010101010110101"; --    -452608   +6695605
      WHEN 2038 => Ti := "111110011011100010000100011001100011010100010000"; --    -411516   +6698256
      WHEN 2039 => Ti := "111110100101100100011000011001100011111001101111"; --    -370408   +6700655
      WHEN 2040 => Ti := "111110101111100110111001011001100100011011010010"; --    -329287   +6702802
      WHEN 2041 => Ti := "111110111001101001100111011001100100111000111000"; --    -288153   +6704696
      WHEN 2042 => Ti := "111111000011101100011111011001100101010010100010"; --    -247009   +6706338
      WHEN 2043 => Ti := "111111001101101111100001011001100101101000001111"; --    -205855   +6707727
      WHEN 2044 => Ti := "111111010111110010101011011001100101111010000000"; --    -164693   +6708864
      WHEN 2045 => Ti := "111111100001110101111011011001100110000111110100"; --    -123525   +6709748
      WHEN 2046 => Ti := "111111101011111001010000011001100110010001101100"; --     -82352   +6710380
      WHEN 2047 => Ti := "111111110101111100100111011001100110010111100111"; --     -41177   +6710759
      WHEN OTHERS => NULL;
    END CASE; 
    T <= Ti; 
  END PROCESS; 
END ARCHITECTURE arch_rom; 



-----------------------------------------------------------
LIBRARY IEEE; 
  USE IEEE.std_logic_1164.all; 

ENTITY goldvect1 IS 
  PORT ( 
    A : IN integer; 
    T : OUT std_logic_vector(47 DOWNTO 0));
END ENTITY goldvect1; 

ARCHITECTURE arch_rom OF goldvect1 IS 
BEGIN 
  PROCESS (A) 
    VARIABLE Ti  : std_logic_vector(47 DOWNTO 0); 
  BEGIN 
    CASE A IS  
      WHEN    0 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN    1 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN    2 => Ti := "111111111111111111111110011001100110011001100000"; --         -2   +6710880
      WHEN    3 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN    4 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN    5 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN    6 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN    7 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN    8 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN    9 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   10 => Ti := "000000000000000000000000111111111111111111111110"; --         +0         -2
      WHEN   11 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   12 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   13 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   14 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   15 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   16 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   17 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   18 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   19 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   20 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   21 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   22 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   23 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   24 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   25 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   26 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN   27 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   28 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   29 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   30 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   31 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   32 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   33 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   34 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN   35 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   36 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   37 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   38 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   39 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   40 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   41 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   42 => Ti := "000000000000000000000000111111111111111111111110"; --         +0         -2
      WHEN   43 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   44 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   45 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   46 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   47 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   48 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   49 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   50 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   51 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   52 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   53 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   54 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   55 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   56 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   57 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   58 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN   59 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   60 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   61 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   62 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   63 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   64 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   65 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   66 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN   67 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   68 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   69 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   70 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   71 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   72 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   73 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   74 => Ti := "000000000000000000000000111111111111111111111110"; --         +0         -2
      WHEN   75 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   76 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   77 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   78 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   79 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   80 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   81 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   82 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   83 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   84 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   85 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   86 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   87 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   88 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   89 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   90 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN   91 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   92 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   93 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   94 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   95 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   96 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   97 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   98 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN   99 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  100 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  101 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  102 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  103 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  104 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  105 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  106 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  107 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  108 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  109 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  110 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  111 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  112 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  113 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  114 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  115 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  116 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  117 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  118 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  119 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  120 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  121 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  122 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  123 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  124 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  125 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  126 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  127 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  128 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  129 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  130 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  131 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  132 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  133 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  134 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  135 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  136 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  137 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  138 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  139 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  140 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  141 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  142 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  143 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  144 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  145 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  146 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  147 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  148 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  149 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  150 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  151 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  152 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  153 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  154 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  155 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  156 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  157 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  158 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  159 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  160 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  161 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  162 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  163 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  164 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  165 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  166 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  167 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  168 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  169 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  170 => Ti := "111111111111111111111111111111111111111111111111"; --         -1         -1
      WHEN  171 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  172 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  173 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  174 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  175 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  176 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  177 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  178 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  179 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  180 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  181 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  182 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  183 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  184 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  185 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  186 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  187 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  188 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  189 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  190 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  191 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  192 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  193 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  194 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  195 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  196 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  197 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  198 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  199 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  200 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  201 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  202 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  203 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  204 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  205 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  206 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  207 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  208 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  209 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  210 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  211 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  212 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  213 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  214 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  215 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  216 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  217 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  218 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  219 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  220 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  221 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  222 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  223 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  224 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  225 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  226 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  227 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  228 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  229 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  230 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  231 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  232 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  233 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  234 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  235 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  236 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  237 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  238 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  239 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  240 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  241 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  242 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  243 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  244 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  245 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  246 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  247 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  248 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  249 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  250 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  251 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  252 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  253 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  254 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  255 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  256 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  257 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  258 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN  259 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  260 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  261 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  262 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  263 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  264 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  265 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  266 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  267 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  268 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  269 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  270 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  271 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  272 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  273 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  274 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  275 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  276 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  277 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  278 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  279 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  280 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  281 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  282 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  283 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  284 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  285 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  286 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  287 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  288 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  289 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  290 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  291 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  292 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  293 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  294 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  295 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  296 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  297 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  298 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  299 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  300 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  301 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  302 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  303 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  304 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  305 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  306 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  307 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  308 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  309 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  310 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  311 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  312 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  313 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  314 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  315 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  316 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  317 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  318 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  319 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  320 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  321 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  322 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN  323 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  324 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  325 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  326 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  327 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  328 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  329 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  330 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  331 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  332 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  333 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  334 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  335 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  336 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  337 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  338 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  339 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  340 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  341 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  342 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  343 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  344 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  345 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  346 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  347 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  348 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  349 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  350 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  351 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  352 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  353 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  354 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  355 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  356 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  357 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  358 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  359 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  360 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  361 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  362 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  363 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  364 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  365 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  366 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  367 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  368 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  369 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  370 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  371 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  372 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  373 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  374 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  375 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  376 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  377 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  378 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  379 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  380 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  381 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  382 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  383 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  384 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  385 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  386 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  387 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  388 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  389 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  390 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  391 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  392 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  393 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  394 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  395 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  396 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  397 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  398 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  399 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  400 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  401 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  402 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  403 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  404 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  405 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  406 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  407 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  408 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  409 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  410 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  411 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  412 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  413 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  414 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  415 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  416 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  417 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  418 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  419 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  420 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  421 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  422 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  423 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  424 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  425 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  426 => Ti := "111111111111111111111111111111111111111111111111"; --         -1         -1
      WHEN  427 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  428 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  429 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  430 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  431 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  432 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  433 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  434 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  435 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  436 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  437 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  438 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  439 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  440 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  441 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  442 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  443 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  444 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  445 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  446 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  447 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  448 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  449 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  450 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  451 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  452 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  453 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  454 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  455 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  456 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  457 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  458 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  459 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  460 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  461 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  462 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  463 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  464 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  465 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  466 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  467 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  468 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  469 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  470 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  471 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  472 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  473 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  474 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  475 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  476 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  477 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  478 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  479 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  480 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  481 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  482 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  483 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  484 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  485 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  486 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  487 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  488 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  489 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  490 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  491 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  492 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  493 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  494 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  495 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  496 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  497 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  498 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  499 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  500 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  501 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  502 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  503 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  504 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  505 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  506 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  507 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  508 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  509 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  510 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  511 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  512 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  513 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  514 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN  515 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  516 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  517 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  518 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  519 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  520 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  521 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  522 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  523 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  524 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  525 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  526 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  527 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  528 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  529 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  530 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  531 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  532 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  533 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  534 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  535 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  536 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  537 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  538 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  539 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  540 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  541 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  542 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  543 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  544 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  545 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  546 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  547 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  548 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  549 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  550 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  551 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  552 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  553 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  554 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  555 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  556 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  557 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  558 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  559 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  560 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  561 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  562 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  563 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  564 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  565 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  566 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  567 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  568 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  569 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  570 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  571 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  572 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  573 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  574 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  575 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  576 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  577 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  578 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  579 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  580 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  581 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  582 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  583 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  584 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  585 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  586 => Ti := "000000000000000000000001000000000000000000000000"; --         +1         +0
      WHEN  587 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  588 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  589 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  590 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  591 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  592 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  593 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  594 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  595 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  596 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  597 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  598 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  599 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  600 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  601 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  602 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  603 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  604 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  605 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  606 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  607 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  608 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  609 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  610 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  611 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  612 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  613 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  614 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  615 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  616 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  617 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  618 => Ti := "000000000000000000000001000000000000000000000000"; --         +1         +0
      WHEN  619 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  620 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  621 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  622 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  623 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  624 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  625 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  626 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  627 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  628 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  629 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  630 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  631 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  632 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  633 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  634 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  635 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  636 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  637 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  638 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  639 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  640 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  641 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  642 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  643 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  644 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  645 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  646 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  647 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  648 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  649 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  650 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  651 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  652 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  653 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  654 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  655 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  656 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  657 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  658 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  659 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  660 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  661 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  662 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  663 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  664 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  665 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  666 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  667 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  668 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  669 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  670 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  671 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  672 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  673 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  674 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  675 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  676 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  677 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  678 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  679 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  680 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  681 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  682 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  683 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  684 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  685 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  686 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  687 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  688 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  689 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  690 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  691 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  692 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  693 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  694 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  695 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  696 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  697 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  698 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  699 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  700 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  701 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  702 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  703 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  704 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  705 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  706 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  707 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  708 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  709 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  710 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  711 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  712 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  713 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  714 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  715 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  716 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  717 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  718 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  719 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  720 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  721 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  722 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  723 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  724 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  725 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  726 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  727 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  728 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  729 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  730 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  731 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  732 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  733 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  734 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  735 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  736 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  737 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  738 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  739 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  740 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  741 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  742 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  743 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  744 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  745 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  746 => Ti := "000000000000000000000001000000000000000000000000"; --         +1         +0
      WHEN  747 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  748 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  749 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  750 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  751 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  752 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  753 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  754 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  755 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  756 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  757 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  758 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  759 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  760 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  761 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  762 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  763 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  764 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  765 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  766 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  767 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  768 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  769 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  770 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN  771 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  772 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  773 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  774 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  775 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  776 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  777 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  778 => Ti := "000000000000000000000001111111111111111111111111"; --         +1         -1
      WHEN  779 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  780 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  781 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  782 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  783 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  784 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  785 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  786 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  787 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  788 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  789 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  790 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  791 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  792 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  793 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  794 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  795 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  796 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  797 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  798 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  799 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  800 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  801 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  802 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  803 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  804 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  805 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  806 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  807 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  808 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  809 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  810 => Ti := "000000000000000000000001111111111111111111111111"; --         +1         -1
      WHEN  811 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  812 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  813 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  814 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  815 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  816 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  817 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  818 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  819 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  820 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  821 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  822 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  823 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  824 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  825 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  826 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  827 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  828 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  829 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  830 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  831 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  832 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  833 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  834 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN  835 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  836 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  837 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  838 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  839 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  840 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  841 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  842 => Ti := "000000000000000000000001000000000000000000000000"; --         +1         +0
      WHEN  843 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  844 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  845 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  846 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  847 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  848 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  849 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  850 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  851 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  852 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  853 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  854 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  855 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  856 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  857 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  858 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  859 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  860 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  861 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  862 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  863 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  864 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  865 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  866 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  867 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  868 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  869 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  870 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  871 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  872 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  873 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  874 => Ti := "000000000000000000000001000000000000000000000000"; --         +1         +0
      WHEN  875 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  876 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  877 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  878 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  879 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  880 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  881 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  882 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  883 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  884 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  885 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  886 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  887 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  888 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  889 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  890 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  891 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  892 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  893 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  894 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  895 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  896 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  897 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  898 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  899 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  900 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  901 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  902 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  903 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  904 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  905 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  906 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  907 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  908 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  909 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  910 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  911 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  912 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  913 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  914 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  915 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  916 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  917 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  918 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  919 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  920 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  921 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  922 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  923 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  924 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  925 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  926 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  927 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  928 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  929 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  930 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN  931 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  932 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  933 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  934 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  935 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  936 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  937 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  938 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  939 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  940 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  941 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  942 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  943 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  944 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  945 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  946 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  947 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  948 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  949 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  950 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  951 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  952 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  953 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  954 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  955 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  956 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  957 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  958 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  959 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  960 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  961 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  962 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  963 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  964 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  965 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  966 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  967 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  968 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  969 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  970 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  971 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  972 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  973 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  974 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  975 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  976 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  977 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  978 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  979 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  980 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  981 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  982 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  983 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  984 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  985 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  986 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  987 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  988 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  989 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  990 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  991 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  992 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  993 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  994 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  995 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  996 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  997 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  998 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN  999 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1000 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1001 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1002 => Ti := "000000000000000000000001000000000000000000000000"; --         +1         +0
      WHEN 1003 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1004 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1005 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1006 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1007 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1008 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1009 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1010 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1011 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1012 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1013 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1014 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1015 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1016 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1017 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1018 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1019 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1020 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1021 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1022 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1023 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1024 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1025 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1026 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1027 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1028 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1029 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1030 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1031 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1032 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1033 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1034 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1035 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1036 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1037 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1038 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1039 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1040 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1041 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1042 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1043 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1044 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1045 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1046 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1047 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1048 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1049 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1050 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1051 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1052 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1053 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1054 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1055 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1056 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1057 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1058 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1059 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1060 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1061 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1062 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1063 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1064 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1065 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1066 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1067 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1068 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1069 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1070 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1071 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1072 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1073 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1074 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1075 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1076 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1077 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1078 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1079 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1080 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1081 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1082 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1083 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1084 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1085 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1086 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1087 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1088 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1089 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1090 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1091 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1092 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1093 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1094 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1095 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1096 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1097 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1098 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1099 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1100 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1101 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1102 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1103 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1104 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1105 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1106 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1107 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1108 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1109 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1110 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1111 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1112 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1113 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1114 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1115 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1116 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1117 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1118 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1119 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1120 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1121 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1122 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1123 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1124 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1125 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1126 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1127 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1128 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1129 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1130 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1131 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1132 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1133 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1134 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1135 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1136 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1137 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1138 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1139 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1140 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1141 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1142 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1143 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1144 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1145 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1146 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1147 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1148 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1149 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1150 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1151 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1152 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1153 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1154 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1155 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1156 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1157 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1158 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1159 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1160 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1161 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1162 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1163 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1164 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1165 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1166 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1167 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1168 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1169 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1170 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1171 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1172 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1173 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1174 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1175 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1176 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1177 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1178 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1179 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1180 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1181 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1182 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1183 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1184 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1185 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1186 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1187 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1188 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1189 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1190 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1191 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1192 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1193 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1194 => Ti := "111111111111111111111111000000000000000000000001"; --         -1         +1
      WHEN 1195 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1196 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1197 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1198 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1199 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1200 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1201 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1202 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1203 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1204 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1205 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1206 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1207 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1208 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1209 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1210 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1211 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1212 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1213 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1214 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1215 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1216 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1217 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1218 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1219 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1220 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1221 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1222 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1223 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1224 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1225 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1226 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1227 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1228 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1229 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1230 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1231 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1232 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1233 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1234 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1235 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1236 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1237 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1238 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1239 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1240 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1241 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1242 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1243 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1244 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1245 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1246 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1247 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1248 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1249 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1250 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1251 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1252 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1253 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1254 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1255 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1256 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1257 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1258 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1259 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1260 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1261 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1262 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1263 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1264 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1265 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1266 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1267 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1268 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1269 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1270 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1271 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1272 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1273 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1274 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1275 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1276 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1277 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1278 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1279 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1280 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1281 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1282 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1283 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1284 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1285 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1286 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1287 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1288 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1289 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1290 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1291 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1292 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1293 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1294 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1295 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1296 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1297 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1298 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1299 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1300 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1301 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1302 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1303 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1304 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1305 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1306 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1307 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1308 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1309 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1310 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1311 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1312 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1313 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1314 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1315 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1316 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1317 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1318 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1319 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1320 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1321 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1322 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1323 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1324 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1325 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1326 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1327 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1328 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1329 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1330 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1331 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1332 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1333 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1334 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1335 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1336 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1337 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1338 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1339 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1340 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1341 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1342 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1343 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1344 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1345 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1346 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1347 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1348 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1349 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1350 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1351 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1352 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1353 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1354 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1355 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1356 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1357 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1358 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1359 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1360 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1361 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1362 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1363 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1364 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1365 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1366 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1367 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1368 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1369 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1370 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1371 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1372 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1373 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1374 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1375 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1376 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1377 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1378 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1379 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1380 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1381 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1382 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1383 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1384 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1385 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1386 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1387 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1388 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1389 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1390 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1391 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1392 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1393 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1394 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1395 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1396 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1397 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1398 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1399 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1400 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1401 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1402 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1403 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1404 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1405 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1406 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1407 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1408 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1409 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1410 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1411 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1412 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1413 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1414 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1415 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1416 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1417 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1418 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1419 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1420 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1421 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1422 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1423 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1424 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1425 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1426 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1427 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1428 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1429 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1430 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1431 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1432 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1433 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1434 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1435 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1436 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1437 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1438 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1439 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1440 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1441 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1442 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1443 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1444 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1445 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1446 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1447 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1448 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1449 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1450 => Ti := "111111111111111111111111000000000000000000000001"; --         -1         +1
      WHEN 1451 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1452 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1453 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1454 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1455 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1456 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1457 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1458 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1459 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1460 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1461 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1462 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1463 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1464 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1465 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1466 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1467 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1468 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1469 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1470 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1471 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1472 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1473 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1474 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1475 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1476 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1477 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1478 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1479 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1480 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1481 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1482 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1483 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1484 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1485 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1486 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1487 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1488 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1489 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1490 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1491 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1492 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1493 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1494 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1495 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1496 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1497 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1498 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1499 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1500 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1501 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1502 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1503 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1504 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1505 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1506 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1507 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1508 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1509 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1510 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1511 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1512 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1513 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1514 => Ti := "000000000000000000000000000000000000000000000001"; --         +0         +1
      WHEN 1515 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1516 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1517 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1518 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1519 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1520 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1521 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1522 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1523 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1524 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1525 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1526 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1527 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1528 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1529 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1530 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1531 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1532 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1533 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1534 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1535 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1536 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1537 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1538 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1539 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1540 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1541 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1542 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1543 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1544 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1545 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1546 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1547 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1548 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1549 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1550 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1551 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1552 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1553 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1554 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1555 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1556 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1557 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1558 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1559 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1560 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1561 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1562 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1563 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1564 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1565 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1566 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1567 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1568 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1569 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1570 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1571 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1572 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1573 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1574 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1575 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1576 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1577 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1578 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1579 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1580 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1581 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1582 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1583 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1584 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1585 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1586 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1587 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1588 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1589 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1590 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1591 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1592 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1593 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1594 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1595 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1596 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1597 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1598 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1599 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1600 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1601 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1602 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1603 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1604 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1605 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1606 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1607 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1608 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1609 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1610 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1611 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1612 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1613 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1614 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1615 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1616 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1617 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1618 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1619 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1620 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1621 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1622 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1623 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1624 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1625 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1626 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1627 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1628 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1629 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1630 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1631 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1632 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1633 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1634 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1635 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1636 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1637 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1638 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1639 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1640 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1641 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1642 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1643 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1644 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1645 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1646 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1647 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1648 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1649 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1650 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1651 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1652 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1653 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1654 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1655 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1656 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1657 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1658 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1659 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1660 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1661 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1662 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1663 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1664 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1665 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1666 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1667 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1668 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1669 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1670 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1671 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1672 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1673 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1674 => Ti := "111111111111111111111110000000000000000000000000"; --         -2         +0
      WHEN 1675 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1676 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1677 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1678 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1679 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1680 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1681 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1682 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1683 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1684 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1685 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1686 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1687 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1688 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1689 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1690 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1691 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1692 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1693 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1694 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1695 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1696 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1697 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1698 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1699 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1700 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1701 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1702 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1703 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1704 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1705 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1706 => Ti := "111111111111111111111110000000000000000000000000"; --         -2         +0
      WHEN 1707 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1708 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1709 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1710 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1711 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1712 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1713 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1714 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1715 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1716 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1717 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1718 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1719 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1720 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1721 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1722 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1723 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1724 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1725 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1726 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1727 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1728 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1729 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1730 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1731 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1732 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1733 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1734 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1735 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1736 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1737 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1738 => Ti := "111111111111111111111110000000000000000000000000"; --         -2         +0
      WHEN 1739 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1740 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1741 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1742 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1743 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1744 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1745 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1746 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1747 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1748 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1749 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1750 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1751 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1752 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1753 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1754 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1755 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1756 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1757 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1758 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1759 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1760 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1761 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1762 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1763 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1764 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1765 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1766 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1767 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1768 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1769 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1770 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1771 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1772 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1773 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1774 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1775 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1776 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1777 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1778 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1779 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1780 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1781 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1782 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1783 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1784 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1785 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1786 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1787 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1788 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1789 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1790 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1791 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1792 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1793 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1794 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1795 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1796 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1797 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1798 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1799 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1800 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1801 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1802 => Ti := "111111111111111111111111111111111111111111111111"; --         -1         -1
      WHEN 1803 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1804 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1805 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1806 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1807 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1808 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1809 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1810 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1811 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1812 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1813 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1814 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1815 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1816 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1817 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1818 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1819 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1820 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1821 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1822 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1823 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1824 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1825 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1826 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1827 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1828 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1829 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1830 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1831 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1832 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1833 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1834 => Ti := "111111111111111111111111111111111111111111111111"; --         -1         -1
      WHEN 1835 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1836 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1837 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1838 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1839 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1840 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1841 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1842 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1843 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1844 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1845 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1846 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1847 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1848 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1849 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1850 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1851 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1852 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1853 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1854 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1855 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1856 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1857 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1858 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1859 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1860 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1861 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1862 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1863 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1864 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1865 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1866 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1867 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1868 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1869 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1870 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1871 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1872 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1873 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1874 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1875 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1876 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1877 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1878 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1879 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1880 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1881 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1882 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1883 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1884 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1885 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1886 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1887 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1888 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1889 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1890 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1891 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1892 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1893 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1894 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1895 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1896 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1897 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1898 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 1899 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1900 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1901 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1902 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1903 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1904 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1905 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1906 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1907 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1908 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1909 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1910 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1911 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1912 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1913 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1914 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1915 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1916 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1917 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1918 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1919 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1920 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1921 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1922 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1923 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1924 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1925 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1926 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1927 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1928 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1929 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1930 => Ti := "111111111111111111111110000000000000000000000000"; --         -2         +0
      WHEN 1931 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1932 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1933 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1934 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1935 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1936 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1937 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1938 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1939 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1940 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1941 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1942 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1943 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1944 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1945 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1946 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1947 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1948 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1949 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1950 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1951 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1952 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1953 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1954 => Ti := "000000000000000000000000111111111111111111111111"; --         +0         -1
      WHEN 1955 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1956 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1957 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1958 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1959 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1960 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1961 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1962 => Ti := "111111111111111111111110000000000000000000000000"; --         -2         +0
      WHEN 1963 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1964 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1965 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1966 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1967 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1968 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1969 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1970 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1971 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1972 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1973 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1974 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1975 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1976 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1977 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1978 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1979 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1980 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1981 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1982 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1983 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1984 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1985 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1986 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1987 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1988 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1989 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1990 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1991 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1992 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1993 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1994 => Ti := "111111111111111111111110000000000000000000000000"; --         -2         +0
      WHEN 1995 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1996 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1997 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1998 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 1999 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2000 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2001 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2002 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2003 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2004 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2005 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2006 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2007 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2008 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2009 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2010 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2011 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2012 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2013 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2014 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2015 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2016 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2017 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2018 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2019 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2020 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2021 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2022 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2023 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2024 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2025 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2026 => Ti := "111111111111111111111111000000000000000000000000"; --         -1         +0
      WHEN 2027 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2028 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2029 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2030 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2031 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2032 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2033 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2034 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2035 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2036 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2037 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2038 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2039 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2040 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2041 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2042 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2043 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2044 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2045 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2046 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN 2047 => Ti := "000000000000000000000000000000000000000000000000"; --         +0         +0
      WHEN OTHERS => NULL;
    END CASE; 
    T <= Ti; 
  END PROCESS; 
END ARCHITECTURE arch_rom; 



-----------------------------------------------------------
LIBRARY IEEE; 
  USE IEEE.std_logic_1164.all; 

ENTITY testvect2 IS 
  PORT ( 
    A : IN integer; 
    T : OUT std_logic_vector(47 DOWNTO 0));
END ENTITY testvect2; 

ARCHITECTURE arch_rom OF testvect2 IS 
BEGIN 
  PROCESS (A) 
    VARIABLE Ti  : std_logic_vector(47 DOWNTO 0); 
  BEGIN 
    CASE A IS  
      WHEN    0 => Ti := "000001011100001011101001110011010110011010000100"; --    +377577   -3316092
      WHEN    1 => Ti := "000111101101110111100110111000010001000101100000"; --   +2022886   -2027168
      WHEN    2 => Ti := "111111010011000001010001000010010010111001010000"; --    -184239    +601680
      WHEN    3 => Ti := "001001111100110010000010111100010010010011110100"; --   +2608258    -973580
      WHEN    4 => Ti := "000110001000000011110011001000011000100101001000"; --   +1605875   +2197832
      WHEN    5 => Ti := "001001000000001000000101110111110001101000100001"; --   +2359813   -2155999
      WHEN    6 => Ti := "000000001010001011001011000101100000100000110110"; --     +41675   +1443894
      WHEN    7 => Ti := "110011011001010011001101111011000110011100111110"; --   -3304243   -1284290
      WHEN    8 => Ti := "111100010101111001110000110101101010000111101111"; --    -958864   -2711057
      WHEN    9 => Ti := "110111010000100100101001110111000101101110101010"; --   -2291415   -2335830
      WHEN   10 => Ti := "111110011011000000111100001100101000000011100001"; --    -413636   +3309793
      WHEN   11 => Ti := "110011001000011001100000110110010111011110011001"; --   -3373472   -2525287
      WHEN   12 => Ti := "111100101011111001111000110011100010111101010101"; --    -868744   -3264683
      WHEN   13 => Ti := "000001101000101000100001000000111011011111001000"; --    +428577    +243656
      WHEN   14 => Ti := "000010100011100101101010000010101110010110001101"; --    +670058    +714125
      WHEN   15 => Ti := "000011111111001001011010110111100100101110110110"; --   +1045082   -2208842
      WHEN   16 => Ti := "111100000001101100110101111110110110111110011000"; --   -1041611    -299112
      WHEN   17 => Ti := "000010100100011100000100110100110001110100001101"; --    +673540   -2941683
      WHEN   18 => Ti := "000111100011110100010110000111010111110100110000"; --   +1981718   +1932592
      WHEN   19 => Ti := "111010101111011111100011000000101000001011110100"; --   -1378333    +164596
      WHEN   20 => Ti := "000101100111011010000001001001101111101000110101"; --   +1472129   +2554421
      WHEN   21 => Ti := "001010101101100010010100001011110010100110011010"; --   +2807956   +3090842
      WHEN   22 => Ti := "110110101001111110000001000001001000000101100111"; --   -2449535    +295271
      WHEN   23 => Ti := "111001000010010101010100111111001001011110011111"; --   -1825452    -223329
      WHEN   24 => Ti := "111000011000001011011110001001011001001000101101"; --   -1998114   +2462253
      WHEN   25 => Ti := "001000100111000100101111000111010001110100101101"; --   +2257199   +1908013
      WHEN   26 => Ti := "001100100110101111110101001100110101100110110011"; --   +3304437   +3365299
      WHEN   27 => Ti := "111101000011110000011011000010111110010011000110"; --    -771045    +779462
      WHEN   28 => Ti := "111010100111110101111010111010001000100011000000"; --   -1409670   -1537856
      WHEN   29 => Ti := "110011100111101001101100001000110100111011101100"; --   -3245460   +2313964
      WHEN   30 => Ti := "110101011000100000110000111100111100001101101010"; --   -2783184    -801942
      WHEN   31 => Ti := "110100011100110110110011000100101001111101010101"; --   -3027533   +1220437
      WHEN   32 => Ti := "001010100010001011110110110011100010110000100010"; --   +2761462   -3265502
      WHEN   33 => Ti := "111001111111111000111000111010011000011001100000"; --   -1573320   -1472928
      WHEN   34 => Ti := "000100101101010000000100000010010111101001010001"; --   +1233924    +621137
      WHEN   35 => Ti := "000101100111000110110100001000110000110010000100"; --   +1470900   +2296964
      WHEN   36 => Ti := "111000010001001110101000111111101110111011100000"; --   -2026584     -69920
      WHEN   37 => Ti := "111111000000010100010110000110010110111101111110"; --    -260842   +1666942
      WHEN   38 => Ti := "001011010011111100001001111111000010101110011100"; --   +2965257    -250980
      WHEN   39 => Ti := "110101110010001010100000000110011000000111100101"; --   -2678112   +1671653
      WHEN   40 => Ti := "111100110111111101001010000010101001111001011000"; --    -819382    +695896
      WHEN   41 => Ti := "000010100110100010011111000110001000101010101100"; --    +682143   +1608364
      WHEN   42 => Ti := "111100010000110011010101000001111110001111100001"; --    -979755    +517089
      WHEN   43 => Ti := "111000110001100101001110110111001100101011100000"; --   -1894066   -2307360
      WHEN   44 => Ti := "000111100100010001001001111110001100111110001000"; --   +1983561    -471160
      WHEN   45 => Ti := "001100010110110110001001000000100011101000100110"; --   +3239305    +145958
      WHEN   46 => Ti := "111011110110111100110001000110100011110001001111"; --   -1085647   +1719375
      WHEN   47 => Ti := "000011110101101111110000110111101001001110111000"; --   +1006576   -2190408
      WHEN   48 => Ti := "110100101000110110110111111111111010010101001011"; --   -2978377     -23221
      WHEN   49 => Ti := "111111111011110111111001000101001110111010010110"; --     -16903   +1371798
      WHEN   50 => Ti := "001011010100101000111101110111000110000001110111"; --   +2968125   -2334601
      WHEN   51 => Ti := "001010001011110010001000110110111100010101000001"; --   +2669704   -2374335
      WHEN   52 => Ti := "111010110001010010110001000101000011101010010010"; --   -1370959   +1325714
      WHEN   53 => Ti := "110100110100000011101111111110001111010001010110"; --   -2932497    -461738
      WHEN   54 => Ti := "000100100000001001100110001100000100001001101101"; --   +1180262   +3162733
      WHEN   55 => Ti := "001001011110001000010000110111001111011011100001"; --   +2482704   -2296095
      WHEN   56 => Ti := "000001111010011011110101001000010110101011100001"; --    +501493   +2190049
      WHEN   57 => Ti := "110111100100001110010111111000001101111000101100"; --   -2210921   -2040276
      WHEN   58 => Ti := "111111001011011110000001001000001111010101000100"; --    -215167   +2159940
      WHEN   59 => Ti := "111111111010011011000110110111010011001110101111"; --     -22842   -2280529
      WHEN   60 => Ti := "111101011001010011110000000110000011110001000011"; --    -682768   +1588291
      WHEN   61 => Ti := "000001100100101000100000111010011110011100101111"; --    +412192   -1448145
      WHEN   62 => Ti := "000110010111001101011111000100110010001101011000"; --   +1667935   +1254232
      WHEN   63 => Ti := "111111001011100001001110000101110011001101110000"; --    -214962   +1520496
      WHEN   64 => Ti := "111100011011011001110010110110011101111011001111"; --    -936334   -2498865
      WHEN   65 => Ti := "110011111010010000001100001000101011111110110110"; --   -3169268   +2277302
      WHEN   66 => Ti := "000011111111000011000000000000100011011110111111"; --   +1044672    +145343
      WHEN   67 => Ti := "110101101100010000110111111110001110101110001001"; --   -2702281    -463991
      WHEN   68 => Ti := "001010100110011011111000001011100111110110010110"; --   +2778872   +3046806
      WHEN   69 => Ti := "111011110111101001100101000001011000110010100000"; --   -1082779    +363680
      WHEN   70 => Ti := "111100100111001001110111111111011001010001110001"; --    -888201    -158607
      WHEN   71 => Ti := "111011000111111100100000001001000000001000100100"; --   -1278176   +2359844
      WHEN   72 => Ti := "111001111110001111010001111110111111101011001110"; --   -1580079    -263474
      WHEN   73 => Ti := "111010101000101100010100001100011110111101000100"; --   -1406188   +3272516
      WHEN   74 => Ti := "000001100010001110111000000110001111100001001000"; --    +402360   +1636424
      WHEN   75 => Ti := "000110100000001010010110111000010101011111001000"; --   +1704598   -2009144
      WHEN   76 => Ti := "111101001100010011101011001000110011110010000101"; --    -736021   +2309253
      WHEN   77 => Ti := "001001110011010001111111000000001001000101001111"; --   +2569343     +37199
      WHEN   78 => Ti := "001100011110011100100101110100000001010111000111"; --   +3270437   -3140153
      WHEN   79 => Ti := "110100010011100000010110000001111110100010101110"; --   -3065834    +518318
      WHEN   80 => Ti := "110111111110101110100001000000111010111011111011"; --   -2102367    +241403
      WHEN   81 => Ti := "000011000011101100010000001000111001101011101110"; --    +801552   +2333422
      WHEN   82 => Ti := "111000000100111011010111000100001001110110101111"; --   -2076969   +1088943
      WHEN   83 => Ti := "110110001010110100001111001000111000001110111010"; --   -2577137   +2327482
      WHEN   84 => Ti := "000110000010010110111110110110001000011110010011"; --   +1582526   -2586733
      WHEN   85 => Ti := "001011000110101100000100111011010110111101000100"; --   +2910980   -1216700
      WHEN   86 => Ti := "111011100111110011000101111010101001000110011001"; --   -1147707   -1404519
      WHEN   87 => Ti := "000101110001111010000101110110111010001011011001"; --   +1515141   -2383143
      WHEN   88 => Ti := "000101001000110011011100001000101011111000011100"; --   +1346780   +2276892
      WHEN   89 => Ti := "000110001001000011110100000010101011110110001100"; --   +1609972    +703884
      WHEN   90 => Ti := "110110101101011110000011111001110010011100011110"; --   -2435197   -1628386
      WHEN   91 => Ti := "110100100100101101010000110011010111000000011110"; --   -2995376   -3313634
      WHEN   92 => Ti := "001000110101110001100111000111111101011000001011"; --   +2317415   +2086411
      WHEN   93 => Ti := "110101111110001010100100111000101101011000111000"; --   -2628956   -1911240
      WHEN   94 => Ti := "110011011000000110011001000001011110110010100010"; --   -3309159    +388258
      WHEN   95 => Ti := "111110101001011101110100110110001110110001100011"; --    -354444   -2560925
      WHEN   96 => Ti := "000100100101000000000001000110100100110111101001"; --   +1200129   +1723881
      WHEN   97 => Ti := "110100111001110011110001000001001110110010011101"; --   -2908943    +322717
      WHEN   98 => Ti := "111000001011101000001100111110011111111011000010"; --   -2049524    -393534
      WHEN   99 => Ti := "111010011100011111011100000101001001000111000111"; --   -1456164   +1348039
      WHEN  100 => Ti := "111000111101100101010010111110011111110111110110"; --   -1844910    -393738
      WHEN  101 => Ti := "000000101001011000001001000010000111001100011000"; --    +169481    +553752
      WHEN  102 => Ti := "110111000111001110001100000011011010011100110111"; --   -2329716    +894775
      WHEN  103 => Ti := "001011101010101100010010000000001110011000011110"; --   +3058450     +58910
      WHEN  104 => Ti := "001010101100000010010100000101001000010111000111"; --   +2801812   +1344967
      WHEN  105 => Ti := "111011100111001100101011111000001011100101011110"; --   -1150165   -2049698
      WHEN  106 => Ti := "001100011111010110001100110111111000100101010111"; --   +3274124   -2127529
      WHEN  107 => Ti := "001100100011111111110100111111000001111000000010"; --   +3293172    -254462
      WHEN  108 => Ti := "000011000001000101110110110101110100000111110010"; --    +790902   -2670094
      WHEN  109 => Ti := "111110001101111101101010110101101111000001010111"; --    -467094   -2690985
      WHEN  110 => Ti := "110100010000000110101110001011001010101001010111"; --   -3079762   +2927191
      WHEN  111 => Ti := "111010011011111100001111001010001110001100001110"; --   -1458417   +2679566
      WHEN  112 => Ti := "000110101100110111001110111001001000110010101000"; --   +1756622   -1799000
      WHEN  113 => Ti := "111000001011101011011001111101110101010100011001"; --   -2049319    -568039
      WHEN  114 => Ti := "000010011110101000110101000011011001011100110111"; --    +649781    +890679
      WHEN  115 => Ti := "111110111100110111100010111110111000010100110010"; --    -274974    -293582
      WHEN  116 => Ti := "000011010000101111100010000010100111111001010111"; --    +855010    +687703
      WHEN  117 => Ti := "001000001110101110001100001001001100111011110101"; --   +2157452   +2412277
      WHEN  118 => Ti := "000101011101111101001010000011010100000011001110"; --   +1433418    +868558
      WHEN  119 => Ti := "111100100111011001110111000001110011010101110111"; --    -887177    +472439
      WHEN  120 => Ti := "000101111001110011101110111000000010010010001110"; --   +1547502   -2087794
      WHEN  121 => Ti := "001010001011101110111011000001100001111100001010"; --   +2669499    +401162
      WHEN  122 => Ti := "110111110110010100111000111001100010010010110010"; --   -2136776   -1694542
      WHEN  123 => Ti := "000100111001010000001001000010110011001100101001"; --   +1283081    +733993
      WHEN  124 => Ti := "111100000000010110011011000010010010001111101001"; --   -1047141    +599017
      WHEN  125 => Ti := "110101000100011101011011111111111110100001111111"; --   -2865317      -6017
      WHEN  126 => Ti := "000010101011100101101101000110010010000100010110"; --    +702829   +1646870
      WHEN  127 => Ti := "000100101101001001101011000011001100110110011001"; --   +1233515    +839065
      WHEN  128 => Ti := "110110110101000100011111000111111010100100111101"; --   -2404065   +2074941
      WHEN  129 => Ti := "001001001110100001110001000010000100001100010111"; --   +2418801    +541463
      WHEN  130 => Ti := "000010101111111100001001001010101001111100011000"; --    +720649   +2793240
      WHEN  131 => Ti := "110100000111100011011110000101111100101010100111"; --   -3114786   +1559207
      WHEN  132 => Ti := "001100000000110010110100000100011010100000011100"; --   +3148980   +1157148
      WHEN  133 => Ti := "000001100101011000100000111011011000100000010001"; --    +415264   -1210351
      WHEN  134 => Ti := "110111011101101110010101111011001001011100111111"; --   -2237547   -1272001
      WHEN  135 => Ti := "001001010000101011011000110110000110001110010011"; --   +2427608   -2595949
      WHEN  136 => Ti := "000110000100010011110010001001000111000101011001"; --   +1590514   +2388313
      WHEN  137 => Ti := "111011011000011001011001110111010010001000010101"; --   -1210791   -2285035
      WHEN  138 => Ti := "110100111110010000100110110101010110010111100111"; --   -2890714   -2791961
      WHEN  139 => Ti := "001000000000010100100000000011101110100110100101"; --   +2098464    +977317
      WHEN  140 => Ti := "111110011111001101110000000001010001011111010001"; --    -396432    +333777
      WHEN  141 => Ti := "111010101010001111100001111101110010011101111110"; --   -1399839    -579714
      WHEN  142 => Ti := "111111110101111110010001111111001111001011010100"; --     -41071    -199980
      WHEN  143 => Ti := "111011010010000010111101110111001110011110101110"; --   -1236803   -2299986
      WHEN  144 => Ti := "111011000011000010110111000110001101100100010100"; --   -1298249   +1628436
      WHEN  145 => Ti := "001011100100001100001111001000011110111000010111"; --   +3031823   +2223639
      WHEN  146 => Ti := "000101100100101101001100001001101011010101100111"; --   +1461068   +2536807
      WHEN  147 => Ti := "001011001011011111010011111011000000000000001000"; --   +2930643   -1310712
      WHEN  148 => Ti := "110100101100011101010010110110100100110100111000"; --   -2963630   -2470600
      WHEN  149 => Ti := "000000011100010001101011000111011010100001100100"; --    +115819   +1943652
      WHEN  150 => Ti := "001011011111010101110100000010111011001111111000"; --   +3011956    +766968
      WHEN  151 => Ti := "001001011011011110101001110101001010110001001001"; --   +2471849   -2839479
      WHEN  152 => Ti := "111011010000100010111101000100000011101101000111"; --   -1242947   +1063751
      WHEN  153 => Ti := "111111111100010001100000110110000000000100101010"; --     -15264   -2621142
      WHEN  154 => Ti := "111010011100011001000011111001001000011100001111"; --   -1456573   -1800433
      WHEN  155 => Ti := "000001000111110101001000001010110111101111101010"; --    +294216   +2849770
      WHEN  156 => Ti := "110101111100011010100100000100010010010110110011"; --   -2636124   +1123763
      WHEN  157 => Ti := "111100101101111101000110111111111011011000011000"; --    -860346     -18920
      WHEN  158 => Ti := "000111010100101010101010000000000010011000011001"; --   +1919658      +9753
      WHEN  159 => Ti := "111100110011010000010101000000010110110010001000"; --    -838635     +93320
      WHEN  160 => Ti := "000000101000101011010110000100111011111010001111"; --    +166614   +1293967
      WHEN  161 => Ti := "111101001000010000011101000010110101101111110110"; --    -752611    +744438
      WHEN  162 => Ti := "000101001000100110101000110011011110000000100000"; --   +1345960   -3284960
      WHEN  163 => Ti := "000010111101101001000001110101111001001110001110"; --    +776769   -2649202
      WHEN  164 => Ti := "111111100110000100100100001001011010110010010100"; --    -106204   +2469012
      WHEN  165 => Ti := "111111101110111011000001000110011100110111100110"; --     -69951   +1691110
      WHEN  166 => Ti := "000111000111100100001011111101000011001010100000"; --   +1865995    -773472
      WHEN  167 => Ti := "111100001001110110011111000001011110001000111100"; --   -1008225    +385596
      WHEN  168 => Ti := "000011001010011001000110001011110010010011001101"; --    +828998   +3089613
      WHEN  169 => Ti := "111100100101111101000011110111110101101011110000"; --    -893117   -2139408
      WHEN  170 => Ti := "000110000010100110111110110110101100000001101110"; --   +1583550   -2441106
      WHEN  171 => Ti := "000010101011011111010100001011101011101111111101"; --    +702420   +3062781
      WHEN  172 => Ti := "111011011101001100101000110100000001111101100001"; --   -1191128   -3137695
      WHEN  173 => Ti := "000011011000000101111110110100101111111101110010"; --    +885118   -2949262
      WHEN  174 => Ti := "001000101100101011001010110110101100000001101110"; --   +2280138   -2441106
      WHEN  175 => Ti := "000010010010101111001011001001011100100010010101"; --    +601035   +2476181
      WHEN  176 => Ti := "001000110111111110011100000101110010110000111101"; --   +2326428   +1518653
      WHEN  177 => Ti := "110110001111111101111000110011101100011010001100"; --   -2556040   -3225972
      WHEN  178 => Ti := "000010110011111100001010000101011100010000110101"; --    +737034   +1426485
      WHEN  179 => Ti := "110100101100110011101100111000111000110101101111"; --   -2962196   -1864337
      WHEN  180 => Ti := "000010111111010101110101110111101001001000011110"; --    +783733   -2190818
      WHEN  181 => Ti := "111011001100000110001000111100000011000011101110"; --   -1261176   -1036050
      WHEN  182 => Ti := "000011111011110010111111111100101110100111001011"; --   +1031359    -857653
      WHEN  183 => Ti := "000111101010110100011000000111110111000100111011"; --   +2010392   +2060603
      WHEN  184 => Ti := "000010101010000010100000000000110011000101011111"; --    +696480    +209247
      WHEN  185 => Ti := "001010000100011000011111000111110000001011010010"; --   +2639391   +2032338
      WHEN  186 => Ti := "000011001001010010101100110111000001101000001111"; --    +824492   -2352625
      WHEN  187 => Ti := "111001100000011011111001111101100111101101111010"; --   -1702151    -623750
      WHEN  188 => Ti := "001000111001111110011100110110110100000100111101"; --   +2334620   -2408131
      WHEN  189 => Ti := "111101111101101101100100110101000000110001000101"; --    -533660   -2880443
      WHEN  190 => Ti := "111010110000000010110000000001111111110010101111"; --   -1376080    +523439
      WHEN  191 => Ti := "111000110010010101001110000001010110010101101100"; --   -1890994    +353644
      WHEN  192 => Ti := "110101110110000000111011111011010010100000001111"; --   -2662341   -1234929
      WHEN  193 => Ti := "110110011101011101111101001000000000010100111111"; --   -2500739   +2098495
      WHEN  194 => Ti := "000111001100000100001101111010100110000110011000"; --   +1884429   -1416808
      WHEN  195 => Ti := "000111001110100100001110001010001111001100001110"; --   +1894670   +2683662
      WHEN  196 => Ti := "000010110000110010100011000110010111000100010111"; --    +724131   +1667351
      WHEN  197 => Ti := "001000111100011000000100111100100100000011111010"; --   +2344452    -900870
      WHEN  198 => Ti := "001001000111101110100001111001001010101111011100"; --   +2390945   -1791012
      WHEN  199 => Ti := "111001011001101000101010111001001100010010101010"; --   -1730006   -1784662
      WHEN  200 => Ti := "001100001110011001010010000001001101000101101001"; --   +3204690    +315753
      WHEN  201 => Ti := "110101000110001010001111110100101100100000111110"; --   -2858353   -2963394
      WHEN  202 => Ti := "111101111100000011111101000000110000000010010001"; --    -540419    +196753
      WHEN  203 => Ti := "111001101000110010010110110101101111011110001010"; --   -1667946   -2689142
      WHEN  204 => Ti := "111000111110001000011111001010001001001000111111"; --   -1842657   +2658879
      WHEN  205 => Ti := "110110001101101101110111110111000100011110101010"; --   -2565257   -2340950
      WHEN  206 => Ti := "110101000100000000101000001011001010110110001011"; --   -2867160   +2928011
      WHEN  207 => Ti := "110100100000111101001110110100100001100000111010"; --   -3010738   -3008454
      WHEN  208 => Ti := "001010011011011111000001111011111011100011101011"; --   +2734017   -1066773
      WHEN  209 => Ti := "111110000101110111001101111101100001011101111000"; --    -500275    -649352
      WHEN  210 => Ti := "001000011100011110010001001011100010101001100000"; --   +2213777   +3025504
      WHEN  211 => Ti := "001000100100100001100001000000111111101011111101"; --   +2246753    +260861
      WHEN  212 => Ti := "111101001100010110111000000101000100101101011111"; --    -735816   +1330015
      WHEN  213 => Ti := "110011000111110110010011111001111100111111101111"; --   -3375725   -1585169
      WHEN  214 => Ti := "001011011101001100001101000000110001100010010010"; --   +3003149    +202898
      WHEN  215 => Ti := "111001001011110010001011111101100001100111011110"; --   -1786741    -648738
      WHEN  216 => Ti := "111001100010110010010011000010010011110010110110"; --   -1692525    +605366
      WHEN  217 => Ti := "001011001101100101101101000100110101000111000000"; --   +2939245   +1266112
      WHEN  218 => Ti := "001001110011011000011000111110011101111011000010"; --   +2569752    -401726
      WHEN  219 => Ti := "001011000110100010011110110011100000000110111011"; --   +2910366   -3276357
      WHEN  220 => Ti := "000111001000110111011000000010101101111111110011"; --   +1871320    +712691
      WHEN  221 => Ti := "110110101010000111101000000010000101001111100100"; --   -2448920    +545764
      WHEN  222 => Ti := "111100110100010011100010111001000000101000111111"; --    -834334   -1832385
      WHEN  223 => Ti := "111101101101100000101011110011011011010110111001"; --    -600021   -3295815
      WHEN  224 => Ti := "000011111010000010111110110101011011000111101001"; --   +1024190   -2772503
      WHEN  225 => Ti := "110100101011000000011111001001001101011011110101"; --   -2969569   +2414325
      WHEN  226 => Ti := "000011111101100010111111001000000101010001110100"; --   +1038527   +2118772
      WHEN  227 => Ti := "000111100011111101111100000101000001010111000100"; --   +1982332   +1316292
      WHEN  228 => Ti := "000100100100001001100111000000111000111111001000"; --   +1196647    +233416
      WHEN  229 => Ti := "000100101010100000000011110110111110010001110100"; --   +1222659   -2366348
      WHEN  230 => Ti := "000110111011000100000110000101111101000001000001"; --   +1814790   +1560641
      WHEN  231 => Ti := "001001010000000100111110110100000111010000110000"; --   +2425150   -3115984
      WHEN  232 => Ti := "000101000110011101000001000011110100011001110100"; --   +1337153   +1001076
      WHEN  233 => Ti := "000001001001001011100010110101100000010111101011"; --    +299746   -2750997
      WHEN  234 => Ti := "110100100001000011101000001011100101011111111011"; --   -3010328   +3037179
      WHEN  235 => Ti := "110110101110100111101010111010010110111001011111"; --   -2430486   -1479073
      WHEN  236 => Ti := "000010111000100101110010001100011101000000010000"; --    +756082   +3264528
      WHEN  237 => Ti := "001010101000001111000110111010110011001100110111"; --   +2786246   -1363145
      WHEN  238 => Ti := "000100110010110000000110111100101110100011111110"; --   +1256454    -857858
      WHEN  239 => Ti := "110111000000001110001010111000111010100101110000"; --   -2358390   -1857168
      WHEN  240 => Ti := "000000010111001000000011111001011110011111100100"; --     +94723   -1710108
      WHEN  241 => Ti := "110101101111000111010010001010011010101111011111"; --   -2690606   +2730975
      WHEN  242 => Ti := "111110010100100000111001001010011011010101111001"; --    -440263   +2733433
      WHEN  243 => Ti := "000111000010001101101111110101010111100111101000"; --   +1844079   -2786840
      WHEN  244 => Ti := "001011111101010010110010110111101101110101010011"; --   +3134642   -2171565
      WHEN  245 => Ti := "001001010010111000001100000111001011100111111000"; --   +2436620   +1882616
      WHEN  246 => Ti := "111110101100111010101001111000101101011111010001"; --    -340311   -1910831
      WHEN  247 => Ti := "000110001110101010001111110011011010100000011111"; --   +1632911   -3299297
      WHEN  248 => Ti := "111101010111110110111100110110001111001110010110"; --    -688708   -2559082
      WHEN  249 => Ti := "001100011011001001010111111011010010001001110101"; --   +3256919   -1236363
      WHEN  250 => Ti := "111001011101110010010010110100010011100100000001"; --   -1713006   -3065599
      WHEN  251 => Ti := "111001010110100101011100111000001010011111000100"; --   -1742500   -2054204
      WHEN  252 => Ti := "000010111001001000111111110111001111111000010101"; --    +758335   -2294251
      WHEN  253 => Ti := "001011000011011100000011001001111111000010100010"; --   +2897667   +2617506
      WHEN  254 => Ti := "000110111110001101101110111000010100111011111011"; --   +1827694   -2011397
      WHEN  255 => Ti := "000011110100110110001001000011110110000110101000"; --   +1002889   +1008040
      WHEN  256 => Ti := "111110101011000001000010001010100101111111100011"; --    -348094   +2777059
      WHEN  257 => Ti := "000100000000111111110100001010111001111001010001"; --   +1052660   +2858577
      WHEN  258 => Ti := "000011010011011001001001110111001011011000010011"; --    +865865   -2312685
      WHEN  259 => Ti := "111101110100010000101101000001111001100010101101"; --    -572371    +497837
      WHEN  260 => Ti := "000000110110011110101000001011011101011111111000"; --    +223144   +3004408
      WHEN  261 => Ti := "000000101111101110100101000010001000010101111111"; --    +195493    +558463
      WHEN  262 => Ti := "111101001011001010000100111001110110101001010011"; --    -740732   -1611181
      WHEN  263 => Ti := "110011111100110000001101111100010010010000100111"; --   -3159027    -973785
      WHEN  264 => Ti := "111000000010101110100011000111101011011000000100"; --   -2085981   +2012676
      WHEN  265 => Ti := "111100111110110011100110110101000111100001001000"; --    -791322   -2852792
      WHEN  266 => Ti := "110100110100111101010110000010011100010010111010"; --   -2928810    +640186
      WHEN  267 => Ti := "110111000000001010111101111000011000001111001001"; --   -2358595   -1997879
      WHEN  268 => Ti := "111110101001001010100111000011110100000110100111"; --    -355673    +999847
      WHEN  269 => Ti := "000100110111010110100010000010110010011111110101"; --   +1275298    +731125
      WHEN  270 => Ti := "000100100010010000000000111110100111011011000101"; --   +1188864    -362811
      WHEN  271 => Ti := "001000011010000100101010111101011110000100010000"; --   +2203946    -663280
      WHEN  272 => Ti := "111000000111110001110001000010011110101100100001"; --   -2065295    +650017
      WHEN  273 => Ti := "001001011100000101000011001011101000000011001001"; --   +2474307   +3047625
      WHEN  274 => Ti := "001100010010101100100001111101010110001010100111"; --   +3222305    -695641
      WHEN  275 => Ti := "001001111100011000011100111000000011111111000010"; --   +2606620   -2080830
      WHEN  276 => Ti := "111110010101000100000110000010000001100101111100"; --    -438010    +530812
      WHEN  277 => Ti := "000101001001101001110101000011011000010000000011"; --   +1350261    +885763
      WHEN  278 => Ti := "111010010100101001000000110100100101101010100010"; --   -1488320   -2991454
      WHEN  279 => Ti := "111101011100101010001011111001111110101100100011"; --    -669045   -1578205
      WHEN  280 => Ti := "000101001100011001110110001010001111010101110100"; --   +1361526   +2684276
      WHEN  281 => Ti := "001001111100111011101001000101111101111010101000"; --   +2608873   +1564328
      WHEN  282 => Ti := "111101001011111010000100111101011001001101110101"; --    -737660    -683147
      WHEN  283 => Ti := "111010111010011001001110001010011101010101111010"; --   -1333682   +2741626
      WHEN  284 => Ti := "000001100111101000100001111101010000010000111110"; --    +424481    -719810
      WHEN  285 => Ti := "000101110010111010000101111100010111101010001111"; --   +1519237    -951665
      WHEN  286 => Ti := "000101110111010011101101000110011001100111100101"; --   +1537261   +1677797
      WHEN  287 => Ti := "110110100101000001001100000110001111111010101110"; --   -2469812   +1638062
      WHEN  288 => Ti := "111001111111011000111000111000011100010101100100"; --   -1575368   -1981084
      WHEN  289 => Ti := "001010010101101000100101000100101111010000100100"; --   +2710053   +1242148
      WHEN  290 => Ti := "000000010000111011001101111100101111000011111111"; --     +69325    -855809
      WHEN  291 => Ti := "001010001111100101010110110110000111100100101101"; --   +2685270   -2590419
      WHEN  292 => Ti := "000000010001011011001101111000100001000101100110"; --     +71373   -1961626
      WHEN  293 => Ti := "111110001111010000110111000100000101010011100001"; --    -461769   +1070305
      WHEN  294 => Ti := "110101010100111010010101000100111011000011110101"; --   -2797931   +1290485
      WHEN  295 => Ti := "110100111100111010001100110101010110101110000001"; --   -2896244   -2790527
      WHEN  296 => Ti := "111100000110100011010001110100000001111010010100"; --   -1021743   -3137900
      WHEN  297 => Ti := "000100110111010000001000111011001011110000001101"; --   +1274888   -1262579
      WHEN  298 => Ti := "111101000111101101010000110110111110001000001110"; --    -754864   -2366962
      WHEN  299 => Ti := "000100010011111100101110110101000011100001000110"; --   +1130286   -2869178
      WHEN  300 => Ti := "111000000110010100111110000101111000001010100101"; --   -2071234   +1540773
      WHEN  301 => Ti := "000010110001100101110000000101000101100000101100"; --    +727408   +1333292
      WHEN  302 => Ti := "000000111100000101000100000100000101011001111010"; --    +246084   +1070714
      WHEN  303 => Ti := "000000111110010101000101110101110101011011000000"; --    +255301   -2664768
      WHEN  304 => Ti := "001011111101100101111111110100100101101010100010"; --   +3135871   -2991454
      WHEN  305 => Ti := "001011110110000010101111111111001100101011010011"; --   +3104943    -210221
      WHEN  306 => Ti := "000000100110101110100010000101111100111101110100"; --    +158626   +1560436
      WHEN  307 => Ti := "000100101111111001101100000100101110011010001010"; --   +1244780   +1238666
      WHEN  308 => Ti := "111100111101100000011001111100110110000100000001"; --    -796647    -827135
      WHEN  309 => Ti := "000111101111100100011010110100100110001101101111"; --   +2029850   -2989201
      WHEN  310 => Ti := "110100100100011010000011110111101010001011101011"; --   -2996605   -2186517
      WHEN  311 => Ti := "000111000110000111010111111011010001001101000010"; --   +1860055   -1240254
      WHEN  312 => Ti := "111011010000001100100011111000110000011111010010"; --   -1244381   -1898542
      WHEN  313 => Ti := "110011001111101111111101111111101110011110101101"; --   -3343363     -71763
      WHEN  314 => Ti := "000000000000110111111010111110100101000100101011"; --      +3578    -372437
      WHEN  315 => Ti := "000110011011100111000111000010110101001100101001"; --   +1685959    +742185
      WHEN  316 => Ti := "111011111101111001100111111101100101100001000110"; --   -1057177    -632762
      WHEN  317 => Ti := "001011001000101111010010001000111001000010000111"; --   +2919378   +2330759
      WHEN  318 => Ti := "001100100010110011000000000011010001101001100111"; --   +3288256    +858727
      WHEN  319 => Ti := "000001011010111110110110110100101011111101110001"; --    +372662   -2965647
      WHEN  320 => Ti := "111100111010011101001011001001011011010010010100"; --    -809141   +2471060
      WHEN  321 => Ti := "111010010010011100001100111011001010011001110010"; --   -1497332   -1268110
      WHEN  322 => Ti := "000010101100011100000111110100000000000111000111"; --    +706311   -3145273
      WHEN  323 => Ti := "110011011111010000000010111101010101010100001101"; --   -3279870    -699123
      WHEN  324 => Ti := "111110101011011010101000110100000111001101100011"; --    -346456   -3116189
      WHEN  325 => Ti := "001010111111101000110101001001010010000101011101"; --   +2882101   +2433373
      WHEN  326 => Ti := "000101101000011010000001111101100110110111100000"; --   +1476225    -627232
      WHEN  327 => Ti := "000111101101010001001100000010111110011100101101"; --   +2020428    +780077
      WHEN  328 => Ti := "000001111011010101011011001001101110101111001111"; --    +505179   +2550735
      WHEN  329 => Ti := "110101000010001101011011000010100011010010111100"; --   -2874533    +668860
      WHEN  330 => Ti := "111110110110000100010011000111100111111110011100"; --    -302829   +1998748
      WHEN  331 => Ti := "000010000110100010010011000010011100000110000110"; --    +551059    +639366
      WHEN  332 => Ti := "000111111001110111101011000001111000111111100000"; --   +2072043    +495584
      WHEN  333 => Ti := "111011110011101100110000000100100010101010000101"; --   -1098960   +1190533
      WHEN  334 => Ti := "111001110110101111001110110011100101000110111101"; --   -1610802   -3255875
      WHEN  335 => Ti := "111000111101000010000101111100000100000000100010"; --   -1847163   -1032158
      WHEN  336 => Ti := "111100100001110110101000000111000011101011000010"; --    -909912   +1850050
      WHEN  337 => Ti := "110110000000001101110010001001100101101000110010"; --   -2620558   +2513458
      WHEN  338 => Ti := "000011000111001111011110000101111001001101110011"; --    +816094   +1545075
      WHEN  339 => Ti := "110111101100101000000001001010001101000101110100"; --   -2176511   +2675060
      WHEN  340 => Ti := "001010000110101011101100000001000001111000110001"; --   +2648812    +269873
      WHEN  341 => Ti := "001011101110001111100000000111010010100001100001"; --   +3072992   +1910881
      WHEN  342 => Ti := "001010000101111011101100111000010111101111001001"; --   +2645740   -1999927
      WHEN  343 => Ti := "001011011010111000111111000111101110111011010010"; --   +2993727   +2027218
      WHEN  344 => Ti := "001001110011100101001011001001000011001000100101"; --   +2570571   +2372133
      WHEN  345 => Ti := "110111110000101000000010000011011010100000000100"; --   -2160126    +894980
      WHEN  346 => Ti := "111001110010111100000000000011000111001100110000"; --   -1626368    +815920
      WHEN  347 => Ti := "000101110000011101010001111001101111000010110111"; --   +1509201   -1642313
      WHEN  348 => Ti := "110111011000110100101101000111011111101011001100"; --   -2257619   +1964748
      WHEN  349 => Ti := "111111010100110001010001000101100110000100000101"; --    -177071   +1466629
      WHEN  350 => Ti := "000111101010010001001011110101011001110111101000"; --   +2008139   -2777624
      WHEN  351 => Ti := "110110001100111101110111001001001101110101011100"; --   -2568329   +2415964
      WHEN  352 => Ti := "000001101100001000100010111011001100001001110011"; --    +442914   -1260941
      WHEN  353 => Ti := "000110100001010111001010111111011011010100111111"; --   +1709514    -150209
      WHEN  354 => Ti := "000101101001001101001110111000001110101111000110"; --   +1479502   -2036794
      WHEN  355 => Ti := "110011011001111001100111001100110010101101001011"; --   -3301785   +3353419
      WHEN  356 => Ti := "000100101110000000000101000011111001100000010000"; --   +1236997   +1021968
      WHEN  357 => Ti := "110100110110111010001010110111110001101011101110"; --   -2920822   -2155794
      WHEN  358 => Ti := "000100010101011001100010111010010110111001011111"; --   +1136226   -1479073
      WHEN  359 => Ti := "000001010000110101001011001000110010111011101011"; --    +331083   +2305771
      WHEN  360 => Ti := "000110111101111101101110111100110100100111001101"; --   +1826670    -833075
      WHEN  361 => Ti := "000011010110011111100100111001010001010101111000"; --    +878564   -1763976
      WHEN  362 => Ti := "111000001111111110101000111001001111111100010001"; --   -2031704   -1769711
      WHEN  363 => Ti := "111010001110011000111101001100001011011001110000"; --   -1513923   +3192432
      WHEN  364 => Ti := "000110101101000111001110110011111001110111000100"; --   +1757646   -3170876
      WHEN  365 => Ti := "110100001101101101000111110111001101001000010100"; --   -3089593   -2305516
      WHEN  366 => Ti := "111011111011111001100110110011100011100000100011"; --   -1065370   -3262429
      WHEN  367 => Ti := "111011110011001001100011000011110011010110100111"; --   -1101213    +996775
      WHEN  368 => Ti := "111101101011001101011101111101111011100111101000"; --    -609443    -542232
      WHEN  369 => Ti := "000000111110000001111000110101101000111010111011"; --    +254072   -2715973
      WHEN  370 => Ti := "111011101010100011000110000101001110000111001001"; --   -1136442   +1368521
      WHEN  371 => Ti := "001001011100011110101001000100001001101101001001"; --   +2475945   +1088329
      WHEN  372 => Ti := "000001100110101110111010000001000001101111001011"; --    +420794    +269259
      WHEN  373 => Ti := "111110111011111010101110110100101100110100001011"; --    -278866   -2962165
      WHEN  374 => Ti := "111101111100000011111101111001111110010110001001"; --    -540419   -1579639
      WHEN  375 => Ti := "111111011110000001010101001001011010111011111010"; --    -139179   +2469626
      WHEN  376 => Ti := "000001011111110101010001110101100011100111101100"; --    +392529   -2737684
      WHEN  377 => Ti := "000110111100010000111010000101011110101101101001"; --   +1819706   +1436521
      WHEN  378 => Ti := "001000110010011000000000001001011100011000101110"; --   +2303488   +2475566
      WHEN  379 => Ti := "001001001001000001101111111010110100011100110111"; --   +2396271   -1358025
      WHEN  380 => Ti := "000110001000011101011010000011110101000011011011"; --   +1607514   +1003739
      WHEN  381 => Ti := "000110100111001101100101001000100010000101001100"; --   +1733477   +2236748
      WHEN  382 => Ti := "001010010001000010001010001001101000111111001100"; --   +2691210   +2527180
      WHEN  383 => Ti := "000000010111111110011101001010101011100010110010"; --     +98205   +2799794
      WHEN  384 => Ti := "110101110001000111010011111110100101100100101011"; --   -2682413    -370389
      WHEN  385 => Ti := "001000000101010100100010111100011000011010010000"; --   +2118946    -948592
      WHEN  386 => Ti := "110111010111000001011111111110010001001010111101"; --   -2264993    -453955
      WHEN  387 => Ti := "000011110101111111110000110011010101110000011101"; --   +1007600   -3318755
      WHEN  388 => Ti := "110100101001001010000100000111000111110100101010"; --   -2977148   +1867050
      WHEN  389 => Ti := "111100111000101001111101110101100111100001010100"; --    -816515   -2721708
      WHEN  390 => Ti := "000111101100000001001100000100110100111010001100"; --   +2015308   +1265292
      WHEN  391 => Ti := "110110101010110100011011110111010000110101001000"; --   -2446053   -2290360
      WHEN  392 => Ti := "111011110111111001100101110100100011110000111011"; --   -1081755   -2999237
      WHEN  393 => Ti := "001100000011111001001110110011110010110000101000"; --   +3161678   -3199960
      WHEN  394 => Ti := "110100011000101001111110000011111001100000010000"; --   -3044738   +1021968
      WHEN  395 => Ti := "000011010101001111100011001010101110001100011010"; --    +873443   +2810650
      WHEN  396 => Ti := "110011100011010000000100111110010111101110001100"; --   -3263484    -427124
      WHEN  397 => Ti := "111101000010111101001110111001100001110101111110"; --    -774322   -1696386
      WHEN  398 => Ti := "000111000001110111010110000100000011111101000111"; --   +1842646   +1064775
      WHEN  399 => Ti := "001000001010001110001010110011111001110000101011"; --   +2139018   -3171285
      WHEN  400 => Ti := "000011001111111111100001110110110111001011011000"; --    +851937   -2395432
      WHEN  401 => Ti := "001100001100001100011110000001011010001100000111"; --   +3195678    +369415
      WHEN  402 => Ti := "111000100000101011100001111111001011101011010011"; --   -1963295    -214317
      WHEN  403 => Ti := "000111000010010100001001111011000001000011010101"; --   +1844489   -1306411
      WHEN  404 => Ti := "111111010100001110000100111100000101100110111100"; --    -179324   -1025604
      WHEN  405 => Ti := "110101101000101101101001000010111000100110010001"; --   -2716823    +756113
      WHEN  406 => Ti := "000110010111001010010010001100100001010110101011"; --   +1667730   +3282347
      WHEN  407 => Ti := "111110101100100100001111110111001011100101000110"; --    -341745   -2311866
      WHEN  408 => Ti := "001100100101001100101000000101100010010111010001"; --   +3298088   +1451473
      WHEN  409 => Ti := "000011011100000110000000000111001011000001011110"; --    +901504   +1880158
      WHEN  410 => Ti := "001011001110111100000111000011001110001100110011"; --   +2944775    +844595
      WHEN  411 => Ti := "111010011011100101110110000100111011111010001111"; --   -1459850   +1293967
      WHEN  412 => Ti := "111010011100100010101001000001110101101001000101"; --   -1455959    +481861
      WHEN  413 => Ti := "000101001111111101000101000001010110101000111001"; --   +1376069    +354873
      WHEN  414 => Ti := "000001000000011110101100111001101000001001001110"; --    +264108   -1670578
      WHEN  415 => Ti := "001011011000101100001011111111111011100001111110"; --   +2984715     -18306
      WHEN  416 => Ti := "000110100110011101100101000100011101110110110111"; --   +1730405   +1170871
      WHEN  417 => Ti := "111110011011000111010101000011010001110000000001"; --    -413227    +859137
      WHEN  418 => Ti := "000110000110010011110011000111110001001000000110"; --   +1598707   +2036230
      WHEN  419 => Ti := "111000010000000001110100001100101000101101000111"; --   -2031500   +3312455
      WHEN  420 => Ti := "001010010011011110111110000011011011110000000100"; --   +2701246    +900100
      WHEN  421 => Ti := "001010100001100010010000000010011101001100100000"; --   +2758800    +643872
      WHEN  422 => Ti := "111111100010100111110000000000010000101011101100"; --    -120336     +68332
      WHEN  423 => Ti := "001001110001111011100100111110110101001110010111"; --   +2563812    -306281
      WHEN  424 => Ti := "110111101100011110011010001011011001001100101010"; --   -2177126   +2986794
      WHEN  425 => Ti := "111000001101011000001101111001110001001100011110"; --   -2042355   -1633506
      WHEN  426 => Ti := "001011000110110010011110000110000001010001000010"; --   +2911390   +1578050
      WHEN  427 => Ti := "110100000100100000010000000011010100100011001111"; --   -3127280    +870607
      WHEN  428 => Ti := "110011111001010011011001000011101111001100111111"; --   -3173159    +979775
      WHEN  429 => Ti := "000000111100111000010001000001100011111100001011"; --    +249361    +409355
      WHEN  430 => Ti := "110100100101010011101001111110101111101011001000"; --   -2992919    -329016
      WHEN  431 => Ti := "110110010010000100010010001100110100010110110010"; --   -2547438   +3360178
      WHEN  432 => Ti := "110100010011010000010110000010101100111100100110"; --   -3066858    +708390
      WHEN  433 => Ti := "000011111010100010111110110111101111011110111010"; --   +1026238   -2164806
      WHEN  434 => Ti := "111011000110011100011111111011110101000011101001"; --   -1284321   -1093399
      WHEN  435 => Ti := "111101100001011010001100000100000011010000010011"; --    -649588   +1061907
      WHEN  436 => Ti := "111000101011111000011000111110010000110100100011"; --   -1917416    -455389
      WHEN  437 => Ti := "110111010001011110010000000100101100000110111100"; --   -2287728   +1229244
      WHEN  438 => Ti := "000000000000100001100001000000000011100101001101"; --      +2145     +14669
      WHEN  439 => Ti := "111110001001100111001111000111110111101000001000"; --    -484913   +2062856
      WHEN  440 => Ti := "111011101100111111111010110011011011110000100000"; --   -1126406   -3294176
      WHEN  441 => Ti := "110110010011011010101100111100111100010000110111"; --   -2541908    -801737
      WHEN  442 => Ti := "000101110010010000011110001000011111111011100100"; --   +1516574   +2227940
      WHEN  443 => Ti := "000011011110110110000001001010001000011111011000"; --    +912769   +2656216
      WHEN  444 => Ti := "000000001011101110011000000011111110010110101011"; --     +48024   +1041835
      WHEN  445 => Ti := "000101111000100110111010000110000110111101111000"; --   +1542586   +1601400
      WHEN  446 => Ti := "111110111100000001001000001011110100100011001110"; --    -278456   +3098830
      WHEN  447 => Ti := "110101111000100100001001111100100111100011111100"; --   -2651895    -886532
      WHEN  448 => Ti := "001000000010010100100001001010011110101001000111"; --   +2106657   +2746951
      WHEN  449 => Ti := "110101110010110100000110111110111101100001100111"; --   -2675450    -272281
      WHEN  450 => Ti := "000110100000010000101111001001100100111011111110"; --   +1705007   +2510590
      WHEN  451 => Ti := "111101101011011101011101110100010100011101101000"; --    -608419   -3061912
      WHEN  452 => Ti := "110100101111110000100000001011010010001100100111"; --   -2950112   +2958119
      WHEN  453 => Ti := "111000011010111011011111110111100010011110110101"; --   -1986849   -2218059
      WHEN  454 => Ti := "000010001001010010010100110110010011111011001011"; --    +562324   -2539829
      WHEN  455 => Ti := "000010110101110010100100110110010110010001100101"; --    +744612   -2530203
      WHEN  456 => Ti := "000100101011110011010001000010001010110110000000"; --   +1227985    +568704
      WHEN  457 => Ti := "001010011101000010001110000110000011000001000011"; --   +2740366   +1585219
      WHEN  458 => Ti := "111010101001110101111011000100011101101101010000"; --   -1401477   +1170256
      WHEN  459 => Ti := "111100101100011001111001001000000001101011011001"; --    -866695   +2104025
      WHEN  460 => Ti := "000110110010100000110110001100110110110000011010"; --   +1779766   +3370010
      WHEN  461 => Ti := "110111011000001110010011111000100011010010011010"; --   -2260077   -1952614
      WHEN  462 => Ti := "110111101001101011001100111101010000100000111110"; --   -2188596    -718786
      WHEN  463 => Ti := "111000000001010001101111000010001100010010110100"; --   -2091921    +574644
      WHEN  464 => Ti := "110111111000011110011111001011111001100011001111"; --   -2127969   +3119311
      WHEN  465 => Ti := "111010110010110101111110111101000101110100000111"; --   -1364610    -762617
      WHEN  466 => Ti := "111000000101011011010111110110011010010100110100"; --   -2074921   -2513612
      WHEN  467 => Ti := "000110110000010100000010110100100000000111010011"; --   +1770754   -3014189
      WHEN  468 => Ti := "001001100100010101000110000110110011010100100010"; --   +2508102   +1783074
      WHEN  469 => Ti := "111110011111110100001010110011010111010000011110"; --    -393974   -3312610
      WHEN  470 => Ti := "000111100010000100010101111110001110111110001001"; --   +1974549    -462967
      WHEN  471 => Ti := "111111101011100100100111111111001000010001101011"; --     -83673    -228245
      WHEN  472 => Ti := "111001000111100010001001000110100000001110000001"; --   -1804151   +1704833
      WHEN  473 => Ti := "110101011000101101100011000001101000111100001101"; --   -2782365    +429837
      WHEN  474 => Ti := "001001111001010010000001001010111011000110000101"; --   +2593921   +2863493
      WHEN  475 => Ti := "110100100010011101001111001001010000100101011101"; --   -3004593   +2427229
      WHEN  476 => Ti := "000011001100010101111010111111111000101011100100"; --    +836986     -29980
      WHEN  477 => Ti := "000110010111100011111001000110011100101010110011"; --   +1669369   +1690291
      WHEN  478 => Ti := "001010010011101000100100111001110111011001010011"; --   +2701860   -1608109
      WHEN  479 => Ti := "111000000111110100111110000111100110000001101000"; --   -2065090   +1990760
      WHEN  480 => Ti := "110100010100101101001010000001011110001100001001"; --   -3060918    +385801
      WHEN  481 => Ti := "000111001111110001000001000000101011111011110110"; --   +1899585    +179958
      WHEN  482 => Ti := "110011101000001001101100000101010110000111001100"; --   -3243412   +1401292
      WHEN  483 => Ti := "000001001011011011100011000110000011010100010000"; --    +308963   +1586448
      WHEN  484 => Ti := "001001011011010101000010001010101110010010110011"; --   +2471234   +2811059
      WHEN  485 => Ti := "111010110101001100011001000111101110001000000101"; --   -1354983   +2023941
      WHEN  486 => Ti := "111111010110010100011111111101011011011101110110"; --    -170721    -673930
      WHEN  487 => Ti := "000011101100111111101100110100101010100000111101"; --    +970732   -2971587
      WHEN  488 => Ti := "000110101100000100000001110011010101110000011101"; --   +1753345   -3318755
      WHEN  489 => Ti := "111000101000110001111110000110101011010111101100"; --   -1930114   +1750508
      WHEN  490 => Ti := "110100011111000000011010110111010001111011100010"; --   -3018726   -2285854
      WHEN  491 => Ti := "110011110110010011011000000100011111001010000100"; --   -3185448   +1176196
      WHEN  492 => Ti := "000100111000001100111100111100001011000011110001"; --   +1278780   -1003279
      WHEN  493 => Ti := "111110001011100100000011000111110000001000000110"; --    -476925   +2032134
      WHEN  494 => Ti := "000011010010000101111100001100011100111001110110"; --    +860540   +3264118
      WHEN  495 => Ti := "111111001110010001001111111010111000001100111000"; --    -203697   -1342664
      WHEN  496 => Ti := "110101000010101010001110001001101100111111001110"; --   -2872690   +2543566
      WHEN  497 => Ti := "110110101011011010110101110101111001110100101000"; --   -2443595   -2646744
      WHEN  498 => Ti := "001010100000111000101001110110111110101011011011"; --   +2756137   -2364709
      WHEN  499 => Ti := "111100100101010000001111111011001110001101000001"; --    -895985   -1252543
      WHEN  500 => Ti := "110100001101001001111010001000001001110101000010"; --   -3091846   +2137410
      WHEN  501 => Ti := "111001001001111110111101001000001010011011011100"; --   -1794115   +2139868
      WHEN  502 => Ti := "111001100101000010010100001010010011100010101001"; --   -1683308   +2701481
      WHEN  503 => Ti := "111000010101100101000011111010001101101100101001"; --   -2008765   -1516759
      WHEN  504 => Ti := "001000101011001011001010111001001100001100010000"; --   +2273994   -1785072
      WHEN  505 => Ti := "001001101111001110110000001001101101110010011011"; --   +2552752   +2546843
      WHEN  506 => Ti := "000010100111000010011111001000111100100010001001"; --    +684191   +2345097
      WHEN  507 => Ti := "110111011101000100101110110100010111010111010000"; --   -2240210   -3050032
      WHEN  508 => Ti := "111100000111111001101011111000000001011011110100"; --   -1016213   -2091276
      WHEN  509 => Ti := "110111101111111110011100111110110100011110010111"; --   -2162788    -309353
      WHEN  510 => Ti := "000010111101100101110100001010001101111100001110"; --    +776564   +2678542
      WHEN  511 => Ti := "001010010110100010001100000001010011100010011110"; --   +2713740    +342174
      WHEN  512 => Ti := "000101101101111010000011000000101100101000101001"; --   +1498755    +182825
      WHEN  513 => Ti := "001011110100111111100010001100111001110000011011"; --   +3100642   +3382299
      WHEN  514 => Ti := "001000100001011011000110001001100001101000110000"; --   +2234054   +2497072
      WHEN  515 => Ti := "111100100110001101000011110111000100101011011101"; --    -892093   -2340131
      WHEN  516 => Ti := "110111011000110111111001111010100110010011001011"; --   -2257415   -1415989
      WHEN  517 => Ti := "000110000000001101010111001100001111110110100101"; --   +1573719   +3210661
      WHEN  518 => Ti := "110011110011010110100011000101101010100000111010"; --   -3197533   +1484858
      WHEN  519 => Ti := "000111110100010111101001000011110101010000001110"; --   +2049513   +1004558
      WHEN  520 => Ti := "000111111101010100011111000110001010001010101100"; --   +2086175   +1614508
      WHEN  521 => Ti := "000101011010101001111100110110100000100100110110"; --   +1419900   -2488010
      WHEN  522 => Ti := "000011101001011111101011111100111010111010011101"; --    +956395    -807267
      WHEN  523 => Ti := "001001110010011110110001001010110000010010110100"; --   +2566065   +2819252
      WHEN  524 => Ti := "000110110100000111010001110100001001000011111101"; --   +1786321   -3108611
      WHEN  525 => Ti := "110011001101001001100010111110110011110100110000"; --   -3354014    -312016
      WHEN  526 => Ti := "111101101110011010010001111001001010111100010000"; --    -596335   -1790192
      WHEN  527 => Ti := "001010100010100101011101110111010100111011100011"; --   +2763101   -2273565
      WHEN  528 => Ti := "111001001110101011110010000000001010011000011100"; --   -1774862     +42524
      WHEN  529 => Ti := "001010001110000101010101000110101000100100011110"; --   +2679125   +1739038
      WHEN  530 => Ti := "110011110101010110100100111000110010001000111001"; --   -3189340   -1891783
      WHEN  531 => Ti := "111000110110101110110110000111000011111011000010"; --   -1872970   +1851074
      WHEN  532 => Ti := "000111101010000001001011000001100100010101110001"; --   +2007115    +410993
      WHEN  533 => Ti := "111011100000000110001111001001001000011000100111"; --   -1179249   +2393639
      WHEN  534 => Ti := "001100011001110010111101000001000111011000110011"; --   +3251389    +292403
      WHEN  535 => Ti := "000011100100101001010000001001100100110010011000"; --    +936528   +2509976
      WHEN  536 => Ti := "000111110100100001001111111001001001011111011100"; --   +2050127   -1796132
      WHEN  537 => Ti := "111100011001111001110010111100110100010100000001"; --    -942478    -834303
      WHEN  538 => Ti := "000001011000011011101000110100001101101010011001"; --    +362216   -3089767
      WHEN  539 => Ti := "110110000101000001000000111101100000010001000100"; --   -2600896    -654268
      WHEN  540 => Ti := "001010000001110010000100111011101000110000010111"; --   +2628740   -1143785
      WHEN  541 => Ti := "001011000101001111010000111000011110011111001100"; --   +2905040   -1972276
      WHEN  542 => Ti := "001000110000010111111111110110100001010001101010"; --   +2295295   -2485142
      WHEN  543 => Ti := "111110011010110100001000001010001101000101110100"; --    -414456   +2675060
      WHEN  544 => Ti := "000011010000110010101111111001000000010010100101"; --    +855215   -1833819
      WHEN  545 => Ti := "000010111111001111011011000001101010000010100111"; --    +783323    +434343
      WHEN  546 => Ti := "110011011011110000000001111110001010100001010100"; --   -3294207    -481196
      WHEN  547 => Ti := "110110100101100001001101001001011100001111001000"; --   -2467763   +2474952
      WHEN  548 => Ti := "111010011111001001000100111010001010011111110100"; --   -1445308   -1529868
      WHEN  549 => Ti := "000001011000101011101000000100110001010000100101"; --    +363240   +1250341
      WHEN  550 => Ti := "000010100011101100000100001011110111011001101000"; --    +670468   +3110504
      WHEN  551 => Ti := "111101110101010111000111000111011111111000000000"; --    -567865   +1965568
      WHEN  552 => Ti := "000101111100010110111100001000010001010001111000"; --   +1557948   +2167928
      WHEN  553 => Ti := "000000001111000100110011110110110010110100111101"; --     +61747   -2413251
      WHEN  554 => Ti := "110011001100001100101110110011110101010000101001"; --   -3357906   -3189719
      WHEN  555 => Ti := "111011100011110011000100000110011110011110000001"; --   -1164092   +1697665
      WHEN  556 => Ti := "111110110110001010101100001010011010011111011111"; --    -302420   +2729951
      WHEN  557 => Ti := "110100010011100000010110000110111110100100100110"; --   -3065834   +1829158
      WHEN  558 => Ti := "110011101000010110011111000011011110001100111001"; --   -3242593    +910137
      WHEN  559 => Ti := "001011110100100101111100000100110010100000100101"; --   +3099004   +1255461
      WHEN  560 => Ti := "000101000110001001110100000000001000010101001111"; --   +1335924     +34127
      WHEN  561 => Ti := "001000000100001010111011111010001000000110001101"; --   +2114235   -1539699
      WHEN  562 => Ti := "000010010011010010011000000011110111110110101001"; --    +603288   +1015209
      WHEN  563 => Ti := "001000101000000001100010111010000100010010111111"; --   +2261090   -1555265
      WHEN  564 => Ti := "000110001010100111000001111111000110001011010001"; --   +1616321    -236847
      WHEN  565 => Ti := "110011011000100000000000111100010100011101011011"; --   -3307520    -964773
      WHEN  566 => Ti := "000011000011001111011101111111100001001011011011"; --    +799709    -126245
      WHEN  567 => Ti := "111100110101010011100010111101101010000111100001"; --    -830238    -613919
      WHEN  568 => Ti := "111010011001111111011011110100000001100111000111"; --   -1466405   -3139129
      WHEN  569 => Ti := "001001101000111110101110000010100110010010111101"; --   +2527150    +681149
      WHEN  570 => Ti := "001010110111000101100101111110011000011110001100"; --   +2847077    -424052
      WHEN  571 => Ti := "000000101010010001110000111101000111110111010101"; --    +173168    -754219
      WHEN  572 => Ti := "001011111101000010110010110011100100110110111101"; --   +3133618   -3256899
      WHEN  573 => Ti := "111110001101011101101010001001011101111111001000"; --    -469142   +2482120
      WHEN  574 => Ti := "111011100010010011000011000101001110101101100011"; --   -1170237   +1370979
      WHEN  575 => Ti := "111111110001100111110110000010101111010011000001"; --     -58890    +718017
      WHEN  576 => Ti := "110100000000101001110101000001101001010010100110"; --   -3143051    +431270
      WHEN  577 => Ti := "111000111110100101010011111101000000000100000101"; --   -1840813    -786171
      WHEN  578 => Ti := "001001000001000100111001001011010100001100101000"; --   +2363705   +2966312
      WHEN  579 => Ti := "000010100110010010011111001100000000000011010010"; --    +681119   +3145938
      WHEN  580 => Ti := "110100111110000000100110000010010001001100011100"; --   -2891738    +594716
      WHEN  581 => Ti := "111010110100111111100101111101101111010001001010"; --   -1355803    -592822
      WHEN  582 => Ti := "110101000011111010001110000000000101010010000001"; --   -2867570     +21633
      WHEN  583 => Ti := "111010110011010010110010001001101101101100000001"; --   -1362766   +2546433
      WHEN  584 => Ti := "001010111001010010011001000111010100110111111011"; --   +2856089   +1920507
      WHEN  585 => Ti := "111000100011000001111100000010011000011111101011"; --   -1953668    +624619
      WHEN  586 => Ti := "000001010111011110110100111010011101111111111011"; --    +358324   -1449989
      WHEN  587 => Ti := "111001011010011111000100001001101101000101101000"; --   -1726524   +2543976
      WHEN  588 => Ti := "000101101000001010000001111011000010001100111100"; --   +1475201   -1301700
      WHEN  589 => Ti := "111000111011011000011110001001100000010010010110"; --   -1853922   +2491542
      WHEN  590 => Ti := "111110011100110100001001111000001100110101011111"; --    -406263   -2044577
      WHEN  591 => Ti := "000001101101110010001010001010000111001100001011"; --    +449674   +2650891
      WHEN  592 => Ti := "001100011111011100100101110100000011100000101110"; --   +3274533   -3131346
      WHEN  593 => Ti := "000010110111010010100101110100110101011010101000"; --    +750757   -2926936
      WHEN  594 => Ti := "110111010111000001011111111001111001010110000111"; --   -2264993   -1600121
      WHEN  595 => Ti := "111000111100000010000101110110010010100111111110"; --   -1851259   -2545154
      WHEN  596 => Ti := "001011100101011001000011111111111111001110110011"; --   +3036739      -3149
      WHEN  597 => Ti := "110101000011001101011011110100100101000111010101"; --   -2870437   -2993707
      WHEN  598 => Ti := "111010001011000101101111111011111101100110111001"; --   -1527441   -1058375
      WHEN  599 => Ti := "111111100100100001010111000000100001000101011000"; --    -112553    +135512
      WHEN  600 => Ti := "001010101011111000101101111101110111110111100111"; --   +2801197    -557593
      WHEN  601 => Ti := "111010011111011100010001000010101101001100100110"; --   -1444079    +709414
      WHEN  602 => Ti := "111101010010110110111010111111011111111000001110"; --    -709190    -131570
      WHEN  603 => Ti := "000001000011001110101101001011101011000110010111"; --    +275373   +3060119
      WHEN  604 => Ti := "000111010110011010101010001000101100011000011100"; --   +1926826   +2278940
      WHEN  605 => Ti := "000010001100001000101110000111110101111000001000"; --    +573998   +2055688
      WHEN  606 => Ti := "111011001001111001010100001001100101111111001011"; --   -1270188   +2514891
      WHEN  607 => Ti := "111001110111101111001110001011010111001100101001"; --   -1606706   +2978601
      WHEN  608 => Ti := "000101011010011101001001001011011101111111111000"; --   +1419081   +3006456
      WHEN  609 => Ti := "000110110110011010011110110110100101011110011110"; --   +1795742   -2467938
      WHEN  610 => Ti := "110111100000111110010110111111011011001011011001"; --   -2224234    -150823
      WHEN  611 => Ti := "110100000100111101000100110100000000000011111010"; --   -3125436   -3145478
      WHEN  612 => Ti := "001001000101101000000111111110111101100001100111"; --   +2382343    -272281
      WHEN  613 => Ti := "110011011000011100110011110110110011011000001010"; --   -3307725   -2410998
      WHEN  614 => Ti := "000111111101111010111001111000110000111111010011"; --   +2088633   -1896493
      WHEN  615 => Ti := "000110111110001101101110000111101110100100111000"; --   +1827694   +2025784
      WHEN  616 => Ti := "111010101010001111100001000100001011010011100011"; --   -1399839   +1094883
      WHEN  617 => Ti := "001010100110101000101011000111010100101110010101"; --   +2779691   +1919893
      WHEN  618 => Ti := "111001001110010010001100001000111000001011101101"; --   -1776500   +2327277
      WHEN  619 => Ti := "110011100110011100111000000000000101100101001110"; --   -3250376     +22862
      WHEN  620 => Ti := "110011110011010110100011110101010000011010110010"; --   -3197533   -2816334
      WHEN  621 => Ti := "000101010100110011100000111100011100000000101011"; --   +1395936    -933845
      WHEN  622 => Ti := "110111101000010111111111111101110011110100011000"; --   -2193921    -574184
      WHEN  623 => Ti := "110111101011001000000000111010111100100000000111"; --   -2182656   -1325049
      WHEN  624 => Ti := "110110011101100001001010000110011000110111100101"; --   -2500534   +1674725
      WHEN  625 => Ti := "000000011101111110011111110100110011110001000001"; --    +122783   -2933695
      WHEN  626 => Ti := "000111101010100100011000111100100000010111000110"; --   +2009368    -916026
      WHEN  627 => Ti := "001010000011001011101011110111011000100101001011"; --   +2634475   -2258613
      WHEN  628 => Ti := "110011110000101001101111110110101100010100111011"; --   -3208593   -2439877
      WHEN  629 => Ti := "000111111101001010111001110111111101101000100110"; --   +2085561   -2106842
      WHEN  630 => Ti := "000001100111110101010100111001101100101100011100"; --    +425300   -1651940
      WHEN  631 => Ti := "000000110101011011011011111100001100110000100101"; --    +218843    -996315
      WHEN  632 => Ti := "001001010011011110100110000100010101110011100111"; --   +2439078   +1137895
      WHEN  633 => Ti := "001011001101100101101101001011001100010010111110"; --   +2939245   +2933950
      WHEN  634 => Ti := "110110111011110100100010110110000000101110010001"; --   -2376414   -2618479
      WHEN  635 => Ti := "000111011111111101111011000001100110100101110010"; --   +1965947    +420210
      WHEN  636 => Ti := "110100110111100011110000001010001111000010101000"; --   -2918160   +2683048
      WHEN  637 => Ti := "001000000100010001010101001001101001101000110011"; --   +2114645   +2529843
      WHEN  638 => Ti := "000001000011111011100000111101010000100100001011"; --    +278240    -718581
      WHEN  639 => Ti := "111110100011100111011000000100100001010110111000"; --    -378408   +1185208
      WHEN  640 => Ti := "001011010100011100001001111010100001011001100011"; --   +2967305   -1436061
      WHEN  641 => Ti := "000101101001101010000001001100011101100110101010"; --   +1481345   +3266986
      WHEN  642 => Ti := "111001111111000010011110000010100010111100100010"; --   -1576802    +667426
      WHEN  643 => Ti := "111000000101000100111101110110101100100100111011"; --   -2076355   -2438853
      WHEN  644 => Ti := "111111011111010001010101000010101100010011000000"; --    -134059    +705728
      WHEN  645 => Ti := "111000111001011110110111111100011010100011110111"; --   -1861705    -939785
      WHEN  646 => Ti := "000100101110010000000101111111100100010001110110"; --   +1238021    -113546
      WHEN  647 => Ti := "000100001100011001011111001011100101111001100010"; --   +1099359   +3038818
      WHEN  648 => Ti := "111001000101111011101111001100011110010011011101"; --   -1810705   +3269853
      WHEN  649 => Ti := "111001000011001000100001000000011101110101010111"; --   -1822175    +122199
      WHEN  650 => Ti := "111111011010010111101101001010010011110010101001"; --    -154131   +2702505
      WHEN  651 => Ti := "000000110001011011011001111011101011010000011000"; --    +202457   -1133544
      WHEN  652 => Ti := "111011101000001001011111000001111011100101111010"; --   -1146273    +506234
      WHEN  653 => Ti := "110111010110000001011111111100001110110011110010"; --   -2269089    -987918
      WHEN  654 => Ti := "111000101000000001111101111010101111110011001111"; --   -1933187   -1377073
      WHEN  655 => Ti := "000101111100101101010101001010111100011001010010"; --   +1559381   +2868818
      WHEN  656 => Ti := "000011101010011111101011000111111110101000001011"; --    +960491   +2091531
      WHEN  657 => Ti := "111001111011010010011101000100111001100000101000"; --   -1592163   +1284136
      WHEN  658 => Ti := "110100101010010011101011000110111100110111110010"; --   -2972437   +1822194
      WHEN  659 => Ti := "001001000000010100111000000101110010111101110000"; --   +2360632   +1519472
      WHEN  660 => Ti := "110100001001011101000101111100000100000000100010"; --   -3107003   -1032158
      WHEN  661 => Ti := "110011100010110011010000111111101101111000010011"; --   -3265328     -74221
      WHEN  662 => Ti := "000010110110001100001011001000110001101110111000"; --    +746251   +2300856
      WHEN  663 => Ti := "000010011110011111001111000001001010000101101000"; --    +649167    +303464
      WHEN  664 => Ti := "000110111010011101101101000001111000001001000110"; --   +1812333    +492102
      WHEN  665 => Ti := "000100110110010110100001000011101101000011011000"; --   +1271201    +970968
      WHEN  666 => Ti := "001001001110111110100100000110110001100001010101"; --   +2420644   +1775701
      WHEN  667 => Ti := "111101110110101010010100110111010111001110110001"; --    -562540   -2264143
      WHEN  668 => Ti := "110011100011110110011110000111011100111110011000"; --   -3261026   +1953688
      WHEN  669 => Ti := "110100000101110011011110111110100010100111110111"; --   -3121954    -382473
      WHEN  670 => Ti := "111001111001111100000011000000010001111011101100"; --   -1597693     +73452
      WHEN  671 => Ti := "111001010001111011110100110101000100001101111010"; --   -1761548   -2866310
      WHEN  672 => Ti := "111111111110100100101110001100011101011101000011"; --      -5842   +3266371
      WHEN  673 => Ti := "110100110101000110111100000011000100111001100010"; --   -2928196    +806498
      WHEN  674 => Ti := "001011011110011001000000111100101110100000110010"; --   +3008064    -858062
      WHEN  675 => Ti := "111011101001101100101100001001010101100101011111"; --   -1139924   +2447711
      WHEN  676 => Ti := "111010011011001001000010111001100000101100011000"; --   -1461694   -1701096
      WHEN  677 => Ti := "001100011011010010111101110100100111110111010110"; --   +3257533   -2982442
      WHEN  678 => Ti := "110100110001101010001000110111101110111011101101"; --   -2942328   -2167059
      WHEN  679 => Ti := "111010101101110010110000111000111101000010100100"; --   -1385296   -1847132
      WHEN  680 => Ti := "000011101001001001010001000111011101100111111111"; --    +954961   +1956351
      WHEN  681 => Ti := "111001101111010010011000110101011101011110000011"; --   -1641320   -2762877
      WHEN  682 => Ti := "111000100101001011100011110110110011111110100100"; --   -1944861   -2408540
      WHEN  683 => Ti := "110111100100110100110001000001101110001001000010"; --   -2208463    +451138
      WHEN  684 => Ti := "110101101111111010011111000011100000010110100000"; --   -2687329    +918944
      WHEN  685 => Ti := "000110011100000111001000111110111011110001100110"; --   +1688008    -279450
      WHEN  686 => Ti := "110100011110110011100111111011110111010011101010"; --   -3019545   -1084182
      WHEN  687 => Ti := "000100110010010110100000111010100011001111111101"; --   +1254816   -1428483
      WHEN  688 => Ti := "000001100010101110111001001001101011001100000000"; --    +404409   +2536192
      WHEN  689 => Ti := "110101000101110011110110001001100011011000110001"; --   -2859786   +2504241
      WHEN  690 => Ti := "001100100110101100101000000111101011101000000100"; --   +3304232   +2013700
      WHEN  691 => Ti := "000010110110101111011000000011100100110011010101"; --    +748504    +937173
      WHEN  692 => Ti := "000010001100100101100010000010100010111001010110"; --    +575842    +667222
      WHEN  693 => Ti := "001100000100101001001111111000010010101000101110"; --   +3164751   -2020818
      WHEN  694 => Ti := "110100000110000011011110111001001111101100010001"; --   -3120930   -1770735
      WHEN  695 => Ti := "111001100010110010010011111001011100000010110000"; --   -1692525   -1720144
      WHEN  696 => Ti := "000111010111010001000100111101101110111010110000"; --   +1930308    -594256
      WHEN  697 => Ti := "001010000011011110111000111010010010110011000100"; --   +2635704   -1495868
      WHEN  698 => Ti := "000101101000110110110100111101000010000100000110"; --   +1478068    -777978
      WHEN  699 => Ti := "110100010111100000010111111000100110101100000010"; --   -3049449   -1938686
      WHEN  700 => Ti := "111100000100110000000011000010110010111100101000"; --   -1029117    +732968
      WHEN  701 => Ti := "000100000111011100101001111100100100010000101110"; --   +1079081    -900050
      WHEN  702 => Ti := "111000101111001011100111001100010011100110100110"; --   -1903897   +3226022
      WHEN  703 => Ti := "111011111001001111111111001010010000000101110101"; --   -1076225   +2687349
      WHEN  704 => Ti := "000100000010100011000001001011101110101100110010"; --   +1059009   +3074866
      WHEN  705 => Ti := "111010001111011000111110111000011110110010011001"; --   -1509826   -1971047
      WHEN  706 => Ti := "000000101000011011010110111100011010110000101010"; --    +165590    -938966
      WHEN  707 => Ti := "111000101001001011100100111010110001001001101001"; --   -1928476   -1371543
      WHEN  708 => Ti := "110101101111100111010010110101110111100100100111"; --   -2688558   -2655961
      WHEN  709 => Ti := "001000100111010100101111000101011110100111001111"; --   +2258223   +1436111
      WHEN  710 => Ti := "000111111110111010111001000100100001001101010010"; --   +2092729   +1184594
      WHEN  711 => Ti := "111111100101110100100100110011011101110011101101"; --    -107228   -3285779
      WHEN  712 => Ti := "001010111101010010011010000010110011000011000010"; --   +2872474    +733378
      WHEN  713 => Ti := "000010100001011000110110111010110000100011001111"; --    +661046   -1374001
      WHEN  714 => Ti := "001001011000100001110101000110011100001010110011"; --   +2459765   +1688243
      WHEN  715 => Ti := "001000010000110111110011001010101011000010110010"; --   +2166259   +2797746
      WHEN  716 => Ti := "111010110100010010110010000010110101001001011100"; --   -1358670    +741980
      WHEN  717 => Ti := "110110110110101110000110000111011001010100110000"; --   -2397306   +1938736
      WHEN  718 => Ti := "000100101001110000000011000001001101011100000010"; --   +1219587    +317186
      WHEN  719 => Ti := "001100011100000110001011111101011010111101110101"; --   +3260811    -675979
      WHEN  720 => Ti := "111101100011001010001101110101111011010111110101"; --    -642419   -2640395
      WHEN  721 => Ti := "000100100111000110011100110100000001010011111010"; --   +1208732   -3140358
      WHEN  722 => Ti := "110111010101101011000101111001111100100010111100"; --   -2270523   -1587012
      WHEN  723 => Ti := "110111110110011011010001111001001010111111011100"; --   -2136367   -1789988
      WHEN  724 => Ti := "000110100011011010010111001001011001000101100000"; --   +1717911   +2462048
      WHEN  725 => Ti := "111111011000100001010011110100100010010111010100"; --    -161709   -3004972
      WHEN  726 => Ti := "001011100111101111011101110100110000010111011001"; --   +3046365   -2947623
      WHEN  727 => Ti := "000001011111010010000100110101011111100111101011"; --    +390276   -2754069
      WHEN  728 => Ti := "000001101101000101010110001011111101100000000100"; --    +446806   +3135492
      WHEN  729 => Ti := "111101011110011010001011001001110100000010011101"; --    -661877   +2572445
      WHEN  730 => Ti := "111101100110010000101000111101101000111010101110"; --    -629720    -618834
      WHEN  731 => Ti := "001000000101110100100010000100001011010110110000"; --   +2120994   +1095088
      WHEN  732 => Ti := "111010010000101000111110001011100001000011000110"; --   -1504706   +3018950
      WHEN  733 => Ti := "000010110010011111010110110011011000000000011110"; --    +731094   -3309538
      WHEN  734 => Ti := "000011110011101100100010110100100101010111010101"; --    +998178   -2992683
      WHEN  735 => Ti := "001011011100101100001100111110000111101110000110"; --   +3001100    -492666
      WHEN  736 => Ti := "111000001001111000001100000010110001111100101000"; --   -2056692    +728872
      WHEN  737 => Ti := "111011101110101111111011111101111011010100011011"; --   -1119237    -543461
      WHEN  738 => Ti := "000111101101010100011001000011010001010110011010"; --   +2020633    +857498
      WHEN  739 => Ti := "110101101101001101101011110011011100010011101101"; --   -2698389   -3291923
      WHEN  740 => Ti := "111010000110011000111010111101011010100111011100"; --   -1546694    -677412
      WHEN  741 => Ti := "001000000111010001010110111011011011011001111001"; --   +2126934   -1198471
      WHEN  742 => Ti := "111010111111001100011100001001001010110101011011"; --   -1314020   +2403675
      WHEN  743 => Ti := "000001011101111110110111111000011000001111001001"; --    +384951   -1997879
      WHEN  744 => Ti := "001100011111001111110010111111010100111011010110"; --   +3273714    -176426
      WHEN  745 => Ti := "111100011100100000001100111110011010001110001101"; --    -931828    -416883
      WHEN  746 => Ti := "111100110111010110110000111110000010100001010001"; --    -821840    -513967
      WHEN  747 => Ti := "001001011110111011011101000010001011011001001101"; --   +2485981    +570957
      WHEN  748 => Ti := "111101000101010011101000111011111101001101010010"; --    -764696   -1060014
      WHEN  749 => Ti := "000000000010111110010101001011101010101001100011"; --     +12181   +3058275
      WHEN  750 => Ti := "000010100101011100000101111110000010001110000100"; --    +677637    -515196
      WHEN  751 => Ti := "110101001001110011110111000111001101000100101100"; --   -2843401   +1888556
      WHEN  752 => Ti := "111000010101011011011101110111001100000101000110"; --   -2009379   -2309818
      WHEN  753 => Ti := "111011001000100110000110110101100011011110000110"; --   -1275514   -2738298
      WHEN  754 => Ti := "000011000111100101111000111111011001011011011000"; --    +817528    -157992
      WHEN  755 => Ti := "110101000010101101011011111011110101100110110110"; --   -2872485   -1091146
      WHEN  756 => Ti := "110110101010110001001111000011000011001111111011"; --   -2446257    +799739
      WHEN  757 => Ti := "001000001000011110001010111010100000010011001001"; --   +2131850   -1440567
      WHEN  758 => Ti := "001100011110000110001011111110100011110001011101"; --   +3269003    -377763
      WHEN  759 => Ti := "110101110000100111010010111000111110011000111110"; --   -2684462   -1841602
      WHEN  760 => Ti := "111001110010010010011001000000100110101111000001"; --   -1629031    +158657
      WHEN  761 => Ti := "000001110000111011110001110011100000011010001000"; --    +462577   -3275128
      WHEN  762 => Ti := "110101110000111010011111000111000010111011000001"; --   -2683233   +1846977
      WHEN  763 => Ti := "111100011110000011011010001100001000011001101111"; --    -925478   +3180143
      WHEN  764 => Ti := "000000010111100100110110001010011101100010101101"; --     +96566   +2742445
      WHEN  765 => Ti := "111010110000100101111101111001000001001100001100"; --   -1373827   -1830132
      WHEN  766 => Ti := "111010111101101100011100111111100100010101000010"; --   -1320164    -113342
      WHEN  767 => Ti := "000110100101110000110010111101111011010111101000"; --   +1727538    -543256
      WHEN  768 => Ti := "111100111110010011100110001000110111010101010011"; --    -793370   +2323795
      WHEN  769 => Ti := "000101100011010011100101111110010000110001010110"; --   +1455333    -455594
      WHEN  770 => Ti := "110101010110100000101111000110001000100001000101"; --   -2791377   +1607749
      WHEN  771 => Ti := "000110010010101010010001110101011010010001001111"; --   +1649297   -2775985
      WHEN  772 => Ti := "000011010101110010110000001001000000001000100100"; --    +875696   +2359844
      WHEN  773 => Ti := "111111001011000100011010111100100001100111000110"; --    -216806    -910906
      WHEN  774 => Ti := "111101101001001101011100110101101111000001010111"; --    -617636   -2690985
      WHEN  775 => Ti := "111011110010111100110000111000001000111111000100"; --   -1102032   -2060348
      WHEN  776 => Ti := "111000111000011110110111001010101100111100011001"; --   -1865801   +2805529
      WHEN  777 => Ti := "110110111101100001010110111011010000110011011011"; --   -2369450   -1241893
      WHEN  778 => Ti := "110111101011011011001101111100000011111101010101"; --   -2181427   -1032363
      WHEN  779 => Ti := "111000010010001011011100111010010010011111110111"; --   -2022692   -1497097
      WHEN  780 => Ti := "111011100110000110010001110111101110111011101101"; --   -1154671   -2167059
      WHEN  781 => Ti := "111111110111000111111000110100111111100100010010"; --     -36360   -2885358
      WHEN  782 => Ti := "000111101110101110000000001011111111010110011110"; --   +2026368   +3143070
      WHEN  783 => Ti := "001010011000101011110011111110101111110111111100"; --   +2722547    -328196
      WHEN  784 => Ti := "111111010110010111101011110111111010000101011000"; --    -170517   -2121384
      WHEN  785 => Ti := "000100111010011100111101111111011001111000001011"; --   +1287997    -156149
      WHEN  786 => Ti := "001010111111100010011011111001101011101100011100"; --   +2881691   -1656036
      WHEN  787 => Ti := "111010101011100010101111111010011010111100101101"; --   -1394513   -1462483
      WHEN  788 => Ti := "000111111111101110000110001000010111111011100001"; --   +2096006   +2195169
      WHEN  789 => Ti := "000111010111011101110111000011011100011100111000"; --   +1931127    +902968
      WHEN  790 => Ti := "111001101100010101100100110011100000001010001000"; --   -1653404   -3276152
      WHEN  791 => Ti := "001011011010001100001011111010101110110000000010"; --   +2990859   -1381374
      WHEN  792 => Ti := "000000010000100100110011001001010100100101011110"; --     +67891   +2443614
      WHEN  793 => Ti := "111001100100011111000111000101011011100111001110"; --   -1685561   +1423822
      WHEN  794 => Ti := "111111100101101010111110001010111001011111101011"; --    -107842   +2856939
      WHEN  795 => Ti := "001000001010000111110001110101101101100111110000"; --   +2138609   -2696720
      WHEN  796 => Ti := "111010001111110101110001110101010010000001001100"; --   -1507983   -2809780
      WHEN  797 => Ti := "000011011110101111100111111101001001010100001000"; --    +912359    -748280
      WHEN  798 => Ti := "111110000011110100000000000000100000010101011000"; --    -508672    +132440
      WHEN  799 => Ti := "001011111110001111100110110110111010111011011010"; --   +3138534   -2380070
      WHEN  800 => Ti := "110011001001001111111010110101001110100111100100"; --   -3369990   -2823708
      WHEN  801 => Ti := "111101100011010000100111001010101111001111100111"; --    -642009   +2814951
      WHEN  802 => Ti := "110111110100001110011101000110101001111110000101"; --   -2145379   +1744773
      WHEN  803 => Ti := "111101110110000011111011110101111011000001011011"; --    -564997   -2641829
      WHEN  804 => Ti := "000000100000111011010011000100101011001010001001"; --    +134867   +1225353
      WHEN  805 => Ti := "001000011100011110010001001000011010110101001001"; --   +2213777   +2207049
      WHEN  806 => Ti := "111111110011001011000011111010010001001100101010"; --     -52541   -1502422
      WHEN  807 => Ti := "110110110100110111101100001001100110100101100101"; --   -2404884   +2517349
      WHEN  808 => Ti := "000000110010111000001101001100001011000000001001"; --    +208397   +3190793
      WHEN  809 => Ti := "110100101110000110111001111000111101111100001011"; --   -2956871   -1843445
      WHEN  810 => Ti := "111000000100101110100011111000100011101000110100"; --   -2077789   -1951180
      WHEN  811 => Ti := "111000000111101011011000111000010000011011111010"; --   -2065704   -2029830
      WHEN  812 => Ti := "000010001101001011111100001011110100000011001101"; --    +578300   +3096781
      WHEN  813 => Ti := "111010100011000101111000000110001110110111100001"; --   -1429128   +1633761
      WHEN  814 => Ti := "000111001000110100001011000100101110010000100011"; --   +1871115   +1238051
      WHEN  815 => Ti := "001010110001111111001001001010111001111100011110"; --   +2826185   +2858782
      WHEN  816 => Ti := "111001101001000101100011001000111011110010001000"; --   -1666717   +2342024
      WHEN  817 => Ti := "110100100110001010000011110110000001000111110111"; --   -2989437   -2616841
      WHEN  818 => Ti := "110110110011110001010010001010011101001100010011"; --   -2409390   +2741011
      WHEN  819 => Ti := "111100001101101001101101001010001011001001000000"; --    -992659   +2667072
      WHEN  820 => Ti := "111100110001111101000111001011110011111001100111"; --    -843961   +3096167
      WHEN  821 => Ti := "000100100010011001100111111011110011011101001111"; --   +1189479   -1099953
      WHEN  822 => Ti := "111100101111100011100000001010000010100101110000"; --    -853792   +2632048
      WHEN  823 => Ti := "000100010010001001100001111110011010010001011010"; --   +1122913    -416678
      WHEN  824 => Ti := "111111010111110111101100111010001001111111110100"; --    -164372   -1531916
      WHEN  825 => Ti := "000111100010111010101111000000110101001111000110"; --   +1978031    +218054
      WHEN  826 => Ti := "000110000111100111000000000111101001100001101010"; --   +1604032   +2005098
      WHEN  827 => Ti := "001000001101000100100101111111110001110001111011"; --   +2150693     -58245
      WHEN  828 => Ti := "111010001001100010100010000001101000010101110011"; --   -1533790    +427379
      WHEN  829 => Ti := "110100011001011101001011111100001101001101011000"; --   -3041461    -994472
      WHEN  830 => Ti := "000110100010110000110000001010101001011100011000"; --   +1715248   +2791192
      WHEN  831 => Ti := "111010001111011100001011111100110000000111001100"; --   -1509621    -851508
      WHEN  832 => Ti := "111011010100100010111110111000101110011111010010"; --   -1226562   -1906734
      WHEN  833 => Ti := "001001100101010001111001110100100110100000111100"; --   +2511993   -2987972
      WHEN  834 => Ti := "111101010110011010001000111001101100000010110110"; --    -694648   -1654602
      WHEN  835 => Ti := "001001011010111000001111110111000001101110101001"; --   +2469391   -2352215
      WHEN  836 => Ti := "000111000100110000111101000010111000101111110111"; --   +1854525    +756727
      WHEN  837 => Ti := "111110100100110111011001111000010110111000101111"; --    -373287   -2003409
      WHEN  838 => Ti := "111110000110110000110100000110110100100001010110"; --    -496588   +1787990
      WHEN  839 => Ti := "000111100111000001001010000011100111001100111100"; --   +1994826    +947004
      WHEN  840 => Ti := "111011010001011100100011110111110010001011101110"; --   -1239261   -2153746
      WHEN  841 => Ti := "000101001011000110101001001011111110100011010001"; --   +1356201   +3139793
      WHEN  842 => Ti := "001001000110100100111011111000011000000010010110"; --   +2386235   -1998698
      WHEN  843 => Ti := "000110000010100000100100110100100001110111010011"; --   +1583140   -3007021
      WHEN  844 => Ti := "110110010111000111100001110100001111011010011001"; --   -2526751   -3082599
      WHEN  845 => Ti := "000001001010010101001001110101011011010100011100"; --    +304457   -2771684
      WHEN  846 => Ti := "000000101010000100111101000001111000100101111001"; --    +172349    +493945
      WHEN  847 => Ti := "110100111111001101011001111000111010111111010110"; --   -2886823   -1855530
      WHEN  848 => Ti := "110100101010010110111000111011000111011100111110"; --   -2972232   -1280194
      WHEN  849 => Ti := "110110011011110100010110111101110110001110000000"; --   -2507498    -564352
      WHEN  850 => Ti := "001000000001010111101101111001110000101111101010"; --   +2102765   -1635350
      WHEN  851 => Ti := "111001111001000010011100000000010101111110111010"; --   -1601380     +90042
      WHEN  852 => Ti := "001010011110011111000010001100100111000110101101"; --   +2746306   +3305901
      WHEN  853 => Ti := "111010010010110010100101110110011011110100110100"; --   -1495899   -2507468
      WHEN  854 => Ti := "111111000100010111100101000101011010101101100111"; --    -244251   +1420135
      WHEN  855 => Ti := "111011110101011100110001111010110111010011010010"; --   -1091791   -1346350
      WHEN  856 => Ti := "000111110001110001001110000000110000101111000100"; --   +2038862    +199620
      WHEN  857 => Ti := "110100101111000011101101000000100011110101011001"; --   -2952979    +146777
      WHEN  858 => Ti := "000001001101001000010111001000100011000001111111"; --    +315927   +2240639
      WHEN  859 => Ti := "000000000011101011001000110101111110001011000011"; --     +15048   -2628925
      WHEN  860 => Ti := "000101100001100011100101001011100011011111111010"; --   +1448165   +3028986
      WHEN  861 => Ti := "111110100100001101110010111111011100111000001100"; --    -375950    -143860
      WHEN  862 => Ti := "000001000100000001111010001010110101111100011100"; --    +278650   +2842396
      WHEN  863 => Ti := "001001101001110001111011111100101010110111001010"; --   +2530427    -873014
      WHEN  864 => Ti := "110110001001100001000010000100001101010011100100"; --   -2582462   +1103076
      WHEN  865 => Ti := "110101111000111101101111000000010011101110111010"; --   -2650257     +80826
      WHEN  866 => Ti := "000001000000001000010010111010011110110011001001"; --    +262674   -1446711
      WHEN  867 => Ti := "111100011101101001110011000111100100111000000001"; --    -927117   +1986049
      WHEN  868 => Ti := "000110000100010110111111001001010010011000101010"; --   +1590719   +2434602
      WHEN  869 => Ti := "111100001110000011010100111111001100011000000110"; --    -991020    -211450
      WHEN  870 => Ti := "000010000000110010010001111110101000101110010011"; --    +527505    -357485
      WHEN  871 => Ti := "000011001100010101111010111101000001011010011111"; --    +836986    -780641
      WHEN  872 => Ti := "111111010111011110000101000001100101111111011000"; --    -166011    +417752
      WHEN  873 => Ti := "110111110001000001101001001000101111001110110111"; --   -2158487   +2290615
      WHEN  874 => Ti := "110101110011110000111010110011100100010000100011"; --   -2671558   -3259357
      WHEN  875 => Ti := "111000101100001000011001110100010110111010011100"; --   -1916391   -3051876
      WHEN  876 => Ti := "111101100001000000100110111001110111101111101101"; --    -651226   -1606675
      WHEN  877 => Ti := "111110010110001010100000000101011011110000110100"; --    -433504   +1424436
      WHEN  878 => Ti := "000000111100001011011101110110101110011000001000"; --    +246493   -2431480
      WHEN  879 => Ti := "000111101010011010110010001001010000001011110110"; --   +2008754   +2425590
      WHEN  880 => Ti := "001010101010011011111010111000111001111111010110"; --   +2795258   -1859626
      WHEN  881 => Ti := "110110101011011010110101111011010101110011011101"; --   -2443595   -1221411
      WHEN  882 => Ti := "110011010001100110010111000010110110101100101010"; --   -3335785    +748330
      WHEN  883 => Ti := "000000110001000001110011001011110010000011001101"; --    +200819   +3088589
      WHEN  884 => Ti := "110011010101000011001011111101001110010000111101"; --   -3321653    -728003
      WHEN  885 => Ti := "001001101011111110101111111001011000110010101110"; --   +2539439   -1733458
      WHEN  886 => Ti := "110110111010110001010101000010011111000110000111"; --   -2380715    +651655
      WHEN  887 => Ti := "000000101101101011011000110011101111011101011010"; --    +187096   -3213478
      WHEN  888 => Ti := "000011101110001111101101001010110010011001001110"; --    +975853   +2827854
      WHEN  889 => Ti := "111101011001010000100011111001000100001001000000"; --    -682973   -1818048
      WHEN  890 => Ti := "110101011111110011111111001100000010110110100000"; --   -2753281   +3157408
      WHEN  891 => Ti := "111111111110000001100001111101100011000100010010"; --      -8095    -642798
      WHEN  892 => Ti := "111011011010110110001101111011111001110000011110"; --   -1200755   -1074146
      WHEN  893 => Ti := "111001011011101000101010000011010101000110011100"; --   -1721814    +872860
      WHEN  894 => Ti := "000000101010111011010111111010101111011100110101"; --    +175831   -1378507
      WHEN  895 => Ti := "111111010000000100011100001010010100110101110110"; --    -196324   +2706806
      WHEN  896 => Ti := "000100010010000011000111111011101110000011100110"; --   +1122503   -1122074
      WHEN  897 => Ti := "000001111011100101011011111111000110101000000100"; --    +506203    -235004
      WHEN  898 => Ti := "001010100111111011111001111101111000101010110100"; --   +2785017    -554316
      WHEN  899 => Ti := "000100000001111001011011110110011010100100110100"; --   +1056347   -2512588
      WHEN  900 => Ti := "111001010110000101011011110111000111111110101011"; --   -1744549   -2326613
      WHEN  901 => Ti := "110101100111111010011100110110001011001011001000"; --   -2720100   -2575672
      WHEN  902 => Ti := "001000001010110111110001000100111110000111000011"; --   +2141681   +1302979
      WHEN  903 => Ti := "111110101000001101110100111111111000011011100100"; --    -359564     -31004
      WHEN  904 => Ti := "111101101110011101011110000100000011000000010011"; --    -596130   +1060883
      WHEN  905 => Ti := "110101100011010100000001000011101100110110100101"; --   -2738943    +970149
      WHEN  906 => Ti := "111100011100110000001100001000100101010010000000"; --    -930804   +2249856
      WHEN  907 => Ti := "000000010100110100110101001001110010111000110111"; --     +85301   +2567735
      WHEN  908 => Ti := "111101000111011101001111001011111101000011010001"; --    -755889   +3133649
      WHEN  909 => Ti := "000011001001111111011111000101111001011010100110"; --    +827359   +1545894
      WHEN  910 => Ti := "000111110101100001001111111100111001010111001111"; --   +2054223    -813617
      WHEN  911 => Ti := "110100101001100000011110001001001001010010001101"; --   -2975714   +2397325
      WHEN  912 => Ti := "111100010010100000001000000110010110101101111110"; --    -972792   +1665918
      WHEN  913 => Ti := "000111111110100111101100111001010110011001000111"; --   +2091500   -1743289
      WHEN  914 => Ti := "111010000001100101101100000111011000011110010110"; --   -1566356   +1935254
      WHEN  915 => Ti := "110111011111000001100010000001101111001100001111"; --   -2232222    +455439
      WHEN  916 => Ti := "000110011001010000101101110110011111111011001111"; --   +1676333   -2490673
      WHEN  917 => Ti := "111010001010100101101111111101111010010111101000"; --   -1529489    -547352
      WHEN  918 => Ti := "000000111100011011011101110111101100011110111001"; --    +247517   -2177095
      WHEN  919 => Ti := "111011001010110010111010111001011111101001001010"; --   -1266502   -1705398
      WHEN  920 => Ti := "000011110110111100100011111001000101001001000001"; --   +1011491   -1813951
      WHEN  921 => Ti := "000100001010111100101011000101001100101101100010"; --   +1093419   +1362786
      WHEN  922 => Ti := "110100011100100011100110000011110010011101000000"; --   -3028762    +993088
      WHEN  923 => Ti := "001011011000111111011000111011110000010000011010"; --   +2985944   -1113062
      WHEN  924 => Ti := "111010111000110010110100111011100001110011100010"; --   -1340236   -1172254
      WHEN  925 => Ti := "111100011100100110100110110111011111011000011010"; --    -931418   -2230758
      WHEN  926 => Ti := "001011100111100010101010111010011001010011000110"; --   +3045546   -1469242
      WHEN  927 => Ti := "111001101100000101100100111001010111011001000111"; --   -1654428   -1739193
      WHEN  928 => Ti := "000110010111100000101100000011010100001001101000"; --   +1669164    +868968
      WHEN  929 => Ti := "111001111100110010011101000010001111010010110101"; --   -1586019    +586933
      WHEN  930 => Ti := "111011101010011001100000000101100011001101101010"; --   -1137056   +1454954
      WHEN  931 => Ti := "110011100100000110011110000101100110011101101100"; --   -3260002   +1468268
      WHEN  932 => Ti := "000011001010001001000110000101010000001101100011"; --    +827974   +1377123
      WHEN  933 => Ti := "000101011100010000010110110110100011011011010001"; --   +1426454   -2476335
      WHEN  934 => Ti := "000000011011001110011110111101000100011101101101"; --    +111518    -768147
      WHEN  935 => Ti := "000010001010101000101110001001011100001111001000"; --    +567854   +2474952
      WHEN  936 => Ti := "110011110011001100111101111111111111101011100110"; --   -3198147      -1306
      WHEN  937 => Ti := "000001001011101000010110000100100001000011101011"; --    +309782   +1183979
      WHEN  938 => Ti := "000001101010111011101111111100010001001010001101"; --    +437999    -978291
      WHEN  939 => Ti := "110011100101110110011110000110111000100111110001"; --   -3252834   +1804785
      WHEN  940 => Ti := "000001000000111011011111110011010101011010000100"; --    +265951   -3320188
      WHEN  941 => Ti := "111010001111001100001010000110011110000100011010"; --   -1510646   +1696026
      WHEN  942 => Ti := "001000011001010001011101000111101001011000000011"; --   +2200669   +2004483
      WHEN  943 => Ti := "111010100110011111100000000101110110010100001011"; --   -1415200   +1533195
      WHEN  944 => Ti := "111101011001010011110000000001000110111100000000"; --    -682768    +290560
      WHEN  945 => Ti := "111100111110110000011001110101111011000111110101"; --    -791527   -2641419
      WHEN  946 => Ti := "000100000111100110010000110101110010110100100101"; --   +1079696   -2675419
      WHEN  947 => Ti := "000100101100110110011110110111011101100010000000"; --   +1232286   -2238336
      WHEN  948 => Ti := "000101111010110011101110000100011111011010000100"; --   +1551598   +1177220
      WHEN  949 => Ti := "000110011000011010010011001010000011101111010110"; --   +1672851   +2636758
      WHEN  950 => Ti := "111001110010110101100110000001111001011111100000"; --   -1626778    +497632
      WHEN  951 => Ti := "111001110110011100000001110110001010111110010100"; --   -1612031   -2576492
      WHEN  952 => Ti := "001100000010010110000001000110000110000111011110"; --   +3155329   +1597918
      WHEN  953 => Ti := "111000100000111000010100111111110011110001111011"; --   -1962476     -50053
      WHEN  954 => Ti := "000010101100111111010100000111110101001000000111"; --    +708564   +2052615
      WHEN  955 => Ti := "111111010111100001010010111100001111011010001100"; --    -165806    -985460
      WHEN  956 => Ti := "111100100101000000001111001100111000011010000001"; --    -897009   +3376769
      WHEN  957 => Ti := "111000101010001110110001001011100101101001100010"; --   -1924175   +3037794
      WHEN  958 => Ti := "000001110000000010001010000011011101000011010010"; --    +458890    +905426
      WHEN  959 => Ti := "001010110100011000110001110111000010110101000011"; --   +2836017   -2347709
      WHEN  960 => Ti := "000011011101001100011010111111000010101011001111"; --    +906010    -251185
      WHEN  961 => Ti := "000011110011001100100010110100100100000100000111"; --    +996130   -2998009
      WHEN  962 => Ti := "110101100100100100000001000110010100110001001010"; --   -2733823   +1657930
      WHEN  963 => Ti := "111000000111110001110001000011111110100110101011"; --   -2065295   +1042859
      WHEN  964 => Ti := "000101110000010110110111111001010100010101111001"; --   +1508791   -1751687
      WHEN  965 => Ti := "000110010100010111000101001100110001111001111110"; --   +1656261   +3350142
      WHEN  966 => Ti := "000001000010000101000110001010001100000010100110"; --    +270662   +2670758
      WHEN  967 => Ti := "001001010000011000001011001010001001100010100101"; --   +2426379   +2660517
      WHEN  968 => Ti := "000101011100010011100011000011000101100110010110"; --   +1426659    +809366
      WHEN  969 => Ti := "110110111001101010111011000110000010001101110110"; --   -2385221   +1581942
      WHEN  970 => Ti := "110110111011000100100001000110101011011010111001"; --   -2379487   +1750713
      WHEN  971 => Ti := "000010101111100101101111111101101011100001001000"; --    +719215    -608184
      WHEN  972 => Ti := "001000010000101011000000000101101010110100000111"; --   +2165440   +1486087
      WHEN  973 => Ti := "110100101001001010000100001010000000001000111100"; --   -2977148   +2622012
      WHEN  974 => Ti := "000010011101110010011011111101011011001010101001"; --    +646299    -675159
      WHEN  975 => Ti := "111110100100010100001100111111110100000101001000"; --    -375540     -48824
      WHEN  976 => Ti := "000001110101000101011001000110110100100100100011"; --    +479577   +1788195
      WHEN  977 => Ti := "000001111100000101011100111011111010011101010001"; --    +508252   -1071279
      WHEN  978 => Ti := "000110001101001101011100111100100010110000101101"; --   +1626972    -906195
      WHEN  979 => Ti := "110101011101011101100101110101011001110100011100"; --   -2762907   -2777828
      WHEN  980 => Ti := "110100001001100110101100001100110110000011100110"; --   -3106388   +3367142
      WHEN  981 => Ti := "110101110010000000111001111101011110010100010000"; --   -2678727    -662256
      WHEN  982 => Ti := "111110000111101101101000111101111100010001001111"; --    -492696    -539569
      WHEN  983 => Ti := "111110100111000001000000111010001110010011000010"; --    -364480   -1514302
      WHEN  984 => Ti := "111001101100111011111110111001000100111111011010"; --   -1650946   -1814566
      WHEN  985 => Ti := "001001111000000101001101000011101111110110100110"; --   +2589005    +982438
      WHEN  986 => Ti := "111110100000111101110001001001110100100010011110"; --    -389263   +2574494
      WHEN  987 => Ti := "111000111100111110111000111101110110111010110011"; --   -1847368    -561485
      WHEN  988 => Ti := "000101111100001101010101001100000000100011010010"; --   +1557333   +3147986
      WHEN  989 => Ti := "000101100001011101001011111100000100010000100010"; --   +1447755   -1031134
      WHEN  990 => Ti := "000010111010111111011010000010110000111111110100"; --    +765914    +724980
      WHEN  991 => Ti := "000100011110111111111111001010001101100010100111"; --   +1175551   +2676903
      WHEN  992 => Ti := "110101110011000000111010111001010110011100010100"; --   -2674630   -1743084
      WHEN  993 => Ti := "000101010101000110101101000000111011011111001000"; --   +1397165    +243656
      WHEN  994 => Ti := "110011011001100000000000000001110110111100010010"; --   -3303424    +487186
      WHEN  995 => Ti := "111110101111111010101010000000011001011110111100"; --    -328022    +104380
      WHEN  996 => Ti := "001001110010011011100101001100001011000110100011"; --   +2565861   +3191203
      WHEN  997 => Ti := "111001010011100010001110000101010011001101100100"; --   -1754994   +1389412
      WHEN  998 => Ti := "111001110101101100000001110101111110000001011100"; --   -1615103   -2629540
      WHEN  999 => Ti := "000010100010111100000100111111010000011000001000"; --    +667396    -195064
      WHEN 1000 => Ti := "111100111001100000010111110100100100110000111011"; --    -813033   -2995141
      WHEN 1001 => Ti := "001100100100001111110100110110010011011110011000"; --   +3294196   -2541672
      WHEN 1002 => Ti := "110100000011101001110110000110010000101101111011"; --   -3130762   +1641339
      WHEN 1003 => Ti := "000100011011010110010111110011011011100011101100"; --   +1160599   -3294996
      WHEN 1004 => Ti := "000101000110100011011011001011110011011100110100"; --   +1337563   +3094324
      WHEN 1005 => Ti := "110110100111111010110100000110100010101010110101"; --   -2457932   +1714869
      WHEN 1006 => Ti := "000010101100101111010100000100101011101101010110"; --    +707540   +1227606
      WHEN 1007 => Ti := "001011111111111100011010000100010010101001111111"; --   +3145498   +1124991
      WHEN 1008 => Ti := "001010001111100010001001110101001000110111100010"; --   +2685065   -2847262
      WHEN 1009 => Ti := "000011000110100010101011001001010111101000101100"; --    +813227   +2456108
      WHEN 1010 => Ti := "000001101111001000100100001010000100111111010111"; --    +455204   +2641879
      WHEN 1011 => Ti := "001010000001001000011101110111001101101110101101"; --   +2626077   -2303059
      WHEN 1012 => Ti := "111001101111100101100101000010000000101100010110"; --   -1640091    +527126
      WHEN 1013 => Ti := "000011000001010010101001110111110011111000100010"; --    +791721   -2146782
      WHEN 1014 => Ti := "000100001010111111111000001000101011011000011100"; --   +1093624   +2274844
      WHEN 1015 => Ti := "111110011111101010100100001001010011001111000100"; --    -394588   +2438084
      WHEN 1016 => Ti := "000011111010010110001011001100011110111101000100"; --   +1025419   +3272516
      WHEN 1017 => Ti := "110100100000001010000001000101011101101010011100"; --   -3014015   +1432220
      WHEN 1018 => Ti := "000110001000100011110011001000001101010101000100"; --   +1607923   +2151748
      WHEN 1019 => Ti := "001000011001011110010000001100010000100000001011"; --   +2201488   +3213323
      WHEN 1020 => Ti := "110110000001100000111111111011010111000011011110"; --   -2615233   -1216290
      WHEN 1021 => Ti := "111010011110110101110111111000100101000101101000"; --   -1446537   -1945240
      WHEN 1022 => Ti := "001000100101001011001000001011100101010011001000"; --   +2249416   +3036360
      WHEN 1023 => Ti := "111000100010100001111011111001101101100110000011"; --   -1955717   -1648253
      WHEN 1024 => Ti := "111110000010110000110010001001011111100101100011"; --    -512974   +2488675
      WHEN 1025 => Ti := "001010110010011111001001111000100101011100000001"; --   +2828233   -1943807
      WHEN 1026 => Ti := "111100111111110000011001000110100110101010110111"; --    -787431   +1731255
      WHEN 1027 => Ti := "000001010010111110110011111100111010010111010000"; --    +339891    -809520
      WHEN 1028 => Ti := "001011000110101100000100000011011101110011010010"; --   +2910980    +908498
      WHEN 1029 => Ti := "000101110110110000100000000110001010101101111001"; --   +1535008   +1616761
      WHEN 1030 => Ti := "000001000110001110101110111101010001010000111111"; --    +287662    -715713
      WHEN 1031 => Ti := "000011000101101100010001001100011010011101000010"; --    +809745   +3254082
      WHEN 1032 => Ti := "111110000001010111001100111011101101010000011001"; --    -518708   -1125351
      WHEN 1033 => Ti := "000100110100100110100001000011011000010000000011"; --   +1264033    +885763
      WHEN 1034 => Ti := "000100000111111001011101111111110111011011100011"; --   +1080925     -35101
      WHEN 1035 => Ti := "110101101100010111010001111010001100000011000001"; --   -2701871   -1523519
      WHEN 1036 => Ti := "110110100101110001001101110100111111001010101011"; --   -2466739   -2886997
      WHEN 1037 => Ti := "110111101000000111111111111110111100001011001101"; --   -2194945    -277811
      WHEN 1038 => Ti := "001000111100100100110111000011110111101001110101"; --   +2345271   +1014389
      WHEN 1039 => Ti := "000111111100010111101100111010001000010110001101"; --   +2082284   -1538675
      WHEN 1040 => Ti := "001010011110111011110101000011010100010000000010"; --   +2748149    +869378
      WHEN 1041 => Ti := "111001100001001111000110110101111011111011000010"; --   -1698874   -2638142
      WHEN 1042 => Ti := "000100111101100011010111000000000010111011100110"; --   +1300695     +12006
      WHEN 1043 => Ti := "110101110100010100000111000101010110000011111111"; --   -2669305   +1401087
      WHEN 1044 => Ti := "111111010110001010111000111100110101110111001110"; --    -171336    -827954
      WHEN 1045 => Ti := "110101100010101101100111001011111011000000000011"; --   -2741401   +3125251
      WHEN 1046 => Ti := "110101011001011010010110111110111101000100110100"; --   -2779498    -274124
      WHEN 1047 => Ti := "111011010110110110001100000000101001100101011011"; --   -1217140    +170331
      WHEN 1048 => Ti := "001000000111000111110000000111100011101000000001"; --   +2126320   +1980929
      WHEN 1049 => Ti := "000001011100110010000011000110001101010001000111"; --    +380035   +1627207
      WHEN 1050 => Ti := "110111110011101110011101110100101001000111010110"; --   -2147427   -2977322
      WHEN 1051 => Ti := "111101111100101101100011001100101011111001111100"; --    -537757   +3325564
      WHEN 1052 => Ti := "000101011110110011100100000011110010100110100111"; --   +1436900    +993703
      WHEN 1053 => Ti := "001000100101111011001000001010011000001111011110"; --   +2252488   +2720734
      WHEN 1054 => Ti := "111111011000000111101100001010110000001001001110"; --    -163348   +2818638
      WHEN 1055 => Ti := "000101101000110000011011111111100110100001110110"; --   +1477659    -104330
      WHEN 1056 => Ti := "111100110101110110101111000110101101110111101101"; --    -827985   +1760749
      WHEN 1057 => Ti := "111010000001101100000101000110011000011010110010"; --   -1565947   +1672882
      WHEN 1058 => Ti := "110011110011111001110000111100100110111101100010"; --   -3195280    -888990
      WHEN 1059 => Ti := "000110011010100011111010001000010111101000010100"; --   +1681658   +2193940
      WHEN 1060 => Ti := "111000110000001110110100111110011100100100101000"; --   -1899596    -407256
      WHEN 1061 => Ti := "111001110100001000110100110101011011011110000011"; --   -1621452   -2771069
      WHEN 1062 => Ti := "000110101001111010011010000011010101100011001111"; --   +1744538    +874703
      WHEN 1063 => Ti := "111001100010000101100000111011101010110000011000"; --   -1695392   -1135592
      WHEN 1064 => Ti := "000110010000101101011101111111101110111110101101"; --   +1641309     -69715
      WHEN 1065 => Ti := "111011111010110011001100000001101101000101110101"; --   -1069876    +446837
      WHEN 1066 => Ti := "001011110001011001000111000101001001010000101110"; --   +3085895   +1348654
      WHEN 1067 => Ti := "111001111111100010011110111101100110100001000111"; --   -1574754    -628665
      WHEN 1068 => Ti := "000010001011010101100001001010000100110010100100"; --    +570721   +2641060
      WHEN 1069 => Ti := "111011111001111001100110000010110110010011000011"; --   -1073562    +746691
      WHEN 1070 => Ti := "001000010000010100100110000111110101011110100001"; --   +2164006   +2054049
      WHEN 1071 => Ti := "111101110110100000101110001000001011101110101010"; --    -563154   +2145194
      WHEN 1072 => Ti := "000011001100111100010100110101011001100001001111"; --    +839444   -2779057
      WHEN 1073 => Ti := "000100101001001001101001001100011110010000010000"; --   +1217129   +3269648
      WHEN 1074 => Ti := "110111101110101011001110000000000110011011101000"; --   -2168114     +26344
      WHEN 1075 => Ti := "111001000111010101010110000001110101110101111000"; --   -1804970    +482680
      WHEN 1076 => Ti := "111010011010001001000010001001011000101111000110"; --   -1465790   +2460614
      WHEN 1077 => Ti := "001000000000001110000111001100101001110000010101"; --   +2098055   +3316757
      WHEN 1078 => Ti := "111011001111111001010110111101100111110111100001"; --   -1245610    -623135
      WHEN 1079 => Ti := "000011110110001100100011111101100001100100010001"; --   +1008419    -648943
      WHEN 1080 => Ti := "001010001001101110111010001011001001100110001010"; --   +2661306   +2922890
      WHEN 1081 => Ti := "000110100100000000110001111010011011010110010100"; --   +1720369   -1460844
      WHEN 1082 => Ti := "001011011001000010100101000000110001101111000101"; --   +2986149    +203717
      WHEN 1083 => Ti := "000011011101011001001101001010110010111001001111"; --    +906829   +2829903
      WHEN 1084 => Ti := "111001110000100101100101110100100010110111010100"; --   -1635995   -3002924
      WHEN 1085 => Ti := "000111010011001101110110111010101101010011001110"; --   +1913718   -1387314
      WHEN 1086 => Ti := "111010010111000010100111111001111011001100100010"; --   -1478489   -1592542
      WHEN 1087 => Ti := "001010011010111111000001111100010100111101011011"; --   +2731969    -962725
      WHEN 1088 => Ti := "111001001111100010001100001000010001011011011111"; --   -1771380   +2168543
      WHEN 1089 => Ti := "111000111001010101010001111011100100001101001001"; --   -1862319   -1162423
      WHEN 1090 => Ti := "111001010010111111000001001011111011010000000011"; --   -1757247   +3126275
      WHEN 1091 => Ti := "000111111101000001010010001011001110000010111111"; --   +2084946   +2941119
      WHEN 1092 => Ti := "000001110010100101011000110101111101110001011100"; --    +469336   -2630564
      WHEN 1093 => Ti := "111100101000110000010001111001001000111001000010"; --    -881647   -1798590
      WHEN 1094 => Ti := "000111001010011010100110111000001101111111000101"; --   +1877670   -2039867
      WHEN 1095 => Ti := "111010111011011100011011001010010001101001000010"; --   -1329381   +2693698
      WHEN 1096 => Ti := "000110010000111101011101110100101101000111011000"; --   +1642333   -2960936
      WHEN 1097 => Ti := "000001010011110101001101000101101110111010100010"; --    +343373   +1502882
      WHEN 1098 => Ti := "111100011100101100111111000001010110001000111001"; --    -931009    +352825
      WHEN 1099 => Ti := "110100110001100110111011110110000111100111111010"; --   -2942533   -2590214
      WHEN 1100 => Ti := "110011101101011001101110000111000111000111110110"; --   -3221906   +1864182
      WHEN 1101 => Ti := "111010111001111100011010111011100000111001111011"; --   -1335526   -1175941
      WHEN 1102 => Ti := "000000011110011110011111110111000001111000001111"; --    +124831   -2351601
      WHEN 1103 => Ti := "000101111110011010001001111011101100100000011001"; --   +1566345   -1128423
      WHEN 1104 => Ti := "000001110110010101011010000010101000111111110001"; --    +484698    +692209
      WHEN 1105 => Ti := "000011111010111001011000001011000001011001010100"; --   +1027672   +2889300
      WHEN 1106 => Ti := "000001111001001011110100000101011111010111001111"; --    +496372   +1439183
      WHEN 1107 => Ti := "111010100011101100010010110101001001111101111100"; --   -1426670   -2842756
      WHEN 1108 => Ti := "000110110001111101101001110011101100010011110011"; --   +1777513   -3226381
      WHEN 1109 => Ti := "000001110110010101011010001100110110101010000000"; --    +484698   +3369600
      WHEN 1110 => Ti := "111111001011001110000001111011001000100000001011"; --    -216191   -1275893
      WHEN 1111 => Ti := "000000001101100100110010110110110001011110100011"; --     +55602   -2418781
      WHEN 1112 => Ti := "000001000101001110101110111000000111001000101001"; --    +283566   -2067927
      WHEN 1113 => Ti := "000000000101111011001001111100111110011101101011"; --     +24265    -792725
      WHEN 1114 => Ti := "000101100001110011100101000100101010001010001000"; --   +1449189   +1221256
      WHEN 1115 => Ti := "000010110001101111010110000101011011110111001110"; --    +728022   +1424846
      WHEN 1116 => Ti := "001011100000101111011011110110011110011110011100"; --   +3017691   -2496612
      WHEN 1117 => Ti := "110100011101000110110011000110000001100001000011"; --   -3026509   +1579075
      WHEN 1118 => Ti := "111111110010000100101001111001001001110101110110"; --     -57047   -1794698
      WHEN 1119 => Ti := "001011111100100010110010110110101111011000001000"; --   +3131570   -2427384
      WHEN 1120 => Ti := "000111000110010111010111111111000000101000000010"; --   +1861079    -259582
      WHEN 1121 => Ti := "000110110110000111010001000010111111011111111010"; --   +1794513    +784378
      WHEN 1122 => Ti := "001000100000000100101100000011000000000110010100"; --   +2228524    +786836
      WHEN 1123 => Ti := "001100100100000011000001111010101101100000000001"; --   +3293377   -1386495
      WHEN 1124 => Ti := "111011101010001111111001001001010001100101011101"; --   -1137671   +2431325
      WHEN 1125 => Ti := "110101110001001101101100110111010110000101001010"; --   -2682004   -2268854
      WHEN 1126 => Ti := "001100000100100110000010001011111110000110011110"; --   +3164546   +3137950
      WHEN 1127 => Ti := "110101111011010000111101000010010001111001001111"; --   -2640835    +597583
      WHEN 1128 => Ti := "111011011110111111110101110101000100100100010100"; --   -1183755   -2864876
      WHEN 1129 => Ti := "111110000010101101100110111101100000110111011110"; --    -513178    -651810
      WHEN 1130 => Ti := "000111100111000001001010000110000111101101111000"; --   +1994826   +1604472
      WHEN 1131 => Ti := "001001011111100001110111000010100110000010111101"; --   +2488439    +680125
      WHEN 1132 => Ti := "001010001111011011101111000001101111111100001111"; --   +2684655    +458511
      WHEN 1133 => Ti := "111000111000010101010000111000100101101111001110"; --   -1866416   -1942578
      WHEN 1134 => Ti := "111110010000101101101011110111111001110101011000"; --    -455829   -2122408
      WHEN 1135 => Ti := "111000100011111011100010111011100001010011100001"; --   -1949982   -1174303
      WHEN 1136 => Ti := "000111000100110100001010001000101100000101001111"; --   +1854730   +2277711
      WHEN 1137 => Ti := "111101001100111101010010001001001111001000101001"; --    -733358   +2421289
      WHEN 1138 => Ti := "001011010011010010100010111110101010100001100000"; --   +2962594    -350112
      WHEN 1139 => Ti := "000111001100100100001101110100100010100000111010"; --   +1886477   -3004358
      WHEN 1140 => Ti := "000000010011111011001110111011000000111001101111"; --     +81614   -1307025
      WHEN 1141 => Ti := "000100001000011001011101111000111110011000111110"; --   +1082973   -1841602
      WHEN 1142 => Ti := "110111011011010100101110111010101111000000000010"; --   -2247378   -1380350
      WHEN 1143 => Ti := "111111000110101010110010001001101001011111001101"; --    -234830   +2529229
      WHEN 1144 => Ti := "001010010110101011110010001000111001010010000111"; --   +2714354   +2331783
      WHEN 1145 => Ti := "110111000101110001011001000010010011010110000011"; --   -2335655    +603523
      WHEN 1146 => Ti := "000100011110001111111111111110101111001011001000"; --   +1172479    -331064
      WHEN 1147 => Ti := "001100001001110110000100001000010000011000010010"; --   +3186052   +2164242
      WHEN 1148 => Ti := "000000001011101011001011001100000010010000000110"; --     +47819   +3154950
      WHEN 1149 => Ti := "110100010011110110110000110101100100100001010011"; --   -3064400   -2733997
      WHEN 1150 => Ti := "001001000101111110100001000010000101100010110001"; --   +2383777    +546993
      WHEN 1151 => Ti := "000010011101010101101000000010011111011100100001"; --    +644456    +653089
      WHEN 1152 => Ti := "111010010000011100001011000010001011100010110011"; --   -1505525    +571571
      WHEN 1153 => Ti := "111100111011000110110001000111100000100001100110"; --    -806479   +1968230
      WHEN 1154 => Ti := "110110000100100111011010001001111000111000111001"; --   -2602534   +2592313
      WHEN 1155 => Ti := "110100011111010110110100001100000110010110100001"; --   -3017292   +3171745
      WHEN 1156 => Ti := "111011110100001001100011111110000001010100011101"; --   -1097117    -518883
      WHEN 1157 => Ti := "110011000011111111111000111100011111110111000110"; --   -3391496    -918074
      WHEN 1158 => Ti := "111000011011011000010010111011011011110110101100"; --   -1985006   -1196628
      WHEN 1159 => Ti := "111111100100110111110001000111010101011011001000"; --    -111119   +1922760
      WHEN 1160 => Ti := "001001110001011000010111110100111000100001000010"; --   +2561559   -2914238
      WHEN 1161 => Ti := "000001100100011000100000111101011111110100010001"; --    +411168    -656111
      WHEN 1162 => Ti := "000101000110011101000001111110101101110111111011"; --   +1337153    -336389
      WHEN 1163 => Ti := "000001111111011011110111000001110111111100010010"; --    +521975    +491282
      WHEN 1164 => Ti := "111000000001001000001000000010110101101001011101"; --   -2092536    +744029
      WHEN 1165 => Ti := "000110111000010000111000111100111011001010011101"; --   +1803320    -806243
      WHEN 1166 => Ti := "000001011101010101010000001010100000100010101110"; --    +382288   +2754734
      WHEN 1167 => Ti := "000111011101101101111010001000000110111110101000"; --   +1956730   +2125736
      WHEN 1168 => Ti := "000110101110101010011011001011100110000011001000"; --   +1763995   +3039432
      WHEN 1169 => Ti := "000011001000111111011111111000010111010101100011"; --    +823263   -2001565
      WHEN 1170 => Ti := "001000100110100001100010000000011110011011110001"; --   +2254946    +124657
      WHEN 1171 => Ti := "000101101011100000011100001000011100010101001001"; --   +1488924   +2213193
      WHEN 1172 => Ti := "000010110110100010100101000100111111111101011101"; --    +747685   +1310557
      WHEN 1173 => Ti := "001001011111111110101010111101011110000100010000"; --   +2490282    -663280
      WHEN 1174 => Ti := "000000101001111000001010001100011110101001110111"; --    +171530   +3271287
      WHEN 1175 => Ti := "000010010111111100000000111001110010111001010010"; --    +622336   -1626542
      WHEN 1176 => Ti := "000011011010101100011001000100101111110011110001"; --    +895769   +1244401
      WHEN 1177 => Ti := "000001011001111110110101001011101010000011001010"; --    +368565   +3055818
      WHEN 1178 => Ti := "000000000100101011001001111010010000111001011101"; --     +19145   -1503651
      WHEN 1179 => Ti := "001001011100000001110110111000100000011000110011"; --   +2474102   -1964493
      WHEN 1180 => Ti := "110110110100111010111001110111101010101011101011"; --   -2404679   -2184469
      WHEN 1181 => Ti := "000100101101110011010001000101110011100000111101"; --   +1236177   +1521725
      WHEN 1182 => Ti := "000010111100001001000000000001100100101100001011"; --    +770624    +412427
      WHEN 1183 => Ti := "001100100111001001011011001100110101000011100110"; --   +3306075   +3363046
      WHEN 1184 => Ti := "000000001010110100110001000010101000011111110001"; --     +44337    +690161
      WHEN 1185 => Ti := "110100001011100110101101000000110000111000101011"; --   -3098195    +200235
      WHEN 1186 => Ti := "001001110111011000011010001000101000101000011011"; --   +2586138   +2263579
      WHEN 1187 => Ti := "111001100101110101100001000001011011010101101110"; --   -1680031    +374126
      WHEN 1188 => Ti := "001010111001111011111111110011011101000110111010"; --   +2858751   -3288646
      WHEN 1189 => Ti := "110101100100010100000001001000001111110101000101"; --   -2734847   +2161989
      WHEN 1190 => Ti := "001000111000110100110101110110101010101110100000"; --   +2329909   -2446432
      WHEN 1191 => Ti := "000110100001110011111101111101000101100111010100"; --   +1711357    -763436
      WHEN 1192 => Ti := "111011010111110010111111110100111111010001000101"; --   -1213249   -2886587
      WHEN 1193 => Ti := "110100111011110011110010110011101110110111000000"; --   -2900750   -3215936
      WHEN 1194 => Ti := "110011001010111111111011111100110010010100000000"; --   -3362821    -842496
      WHEN 1195 => Ti := "000001101110001110111101111001001101011001000100"; --    +451517   -1780156
      WHEN 1196 => Ti := "111100000101111001101010000110011011011010110011"; --   -1024406   +1685171
      WHEN 1197 => Ti := "110101111100110000111101111110100100010100101010"; --   -2634691    -375510
      WHEN 1198 => Ti := "111101000111100011101001001000011111011000010111"; --    -755479   +2225687
      WHEN 1199 => Ti := "001010111011100101100110111011100000011101001000"; --   +2865510   -1177784
      WHEN 1200 => Ti := "000001011101011110110111000010100110110010111101"; --    +382903    +683197
      WHEN 1201 => Ti := "000001111110111000101010001001101010010010011010"; --    +519722   +2532506
      WHEN 1202 => Ti := "111011001111101100100011111001010111101100010100"; --   -1246429   -1737964
      WHEN 1203 => Ti := "000011000011101111011101111001010011111001000110"; --    +801757   -1753530
      WHEN 1204 => Ti := "000011110110100110001010000100000110010000010100"; --   +1010058   +1074196
      WHEN 1205 => Ti := "111111110011010111110110000110110010010100100010"; --     -51722   +1778978
      WHEN 1206 => Ti := "110111100000010111111100000000011010011011101111"; --   -2226692    +108271
      WHEN 1207 => Ti := "111111000100011101111110111110000100010100011110"; --    -243842    -506594
      WHEN 1208 => Ti := "001001101110001000010110001100100001010000010001"; --   +2548246   +3281937
      WHEN 1209 => Ti := "110100111000110011110001110011111000101010010001"; --   -2913039   -3175791
      WHEN 1210 => Ti := "111100111110110000011001110101101100000100100010"; --    -791527   -2703070
      WHEN 1211 => Ti := "001010111000010010011000111011011100000011011111"; --   +2851992   -1195809
      WHEN 1212 => Ti := "000001101100011011101111001000101000001000011011"; --    +444143   +2261531
      WHEN 1213 => Ti := "111101000111011101001111111111111110000101001100"; --    -755889      -7860
      WHEN 1214 => Ti := "000000010111111110011101001010110111010110000011"; --     +98205   +2848131
      WHEN 1215 => Ti := "001001000011011011010011110110001100110111111100"; --   +2373331   -2568708
      WHEN 1216 => Ti := "000110010010010000101010111110000001000111101010"; --   +1647658    -519702
      WHEN 1217 => Ti := "111000110111101011101010001100110011110110110010"; --   -1869078   +3358130
      WHEN 1218 => Ti := "111110111011001101111011110100000101110011111100"; --    -281733   -3121924
      WHEN 1219 => Ti := "111100000111001001101011110110010110010100110010"; --   -1019285   -2529998
      WHEN 1220 => Ti := "001011001011011100000110111100000001110110111010"; --   +2930438   -1040966
      WHEN 1221 => Ti := "001011001000101000111000110011110101110011110110"; --   +2918968   -3187466
      WHEN 1222 => Ti := "000110111001010100000110000111010100010111111011"; --   +1807622   +1918459
      WHEN 1223 => Ti := "000110001110110011110110000111001100010001011111"; --   +1633526   +1885279
      WHEN 1224 => Ti := "110100001000111001111000000011000010100110010101"; --   -3109256    +797077
      WHEN 1225 => Ti := "000001001100100001111101110100101010111010100100"; --    +313469   -2969948
      WHEN 1226 => Ti := "110110011110011101111101000101001011100000101110"; --   -2496643   +1357870
      WHEN 1227 => Ti := "000101101111001101010000111010101001101001100110"; --   +1504080   -1402266
      WHEN 1228 => Ti := "111011111010011100110011111011110001001101001110"; --   -1071309   -1109170
      WHEN 1229 => Ti := "001010010110001011110010000000010111101000100001"; --   +2712306     +96801
      WHEN 1230 => Ti := "001010101100010010010100001011100000001001011111"; --   +2802836   +3015263
      WHEN 1231 => Ti := "000001100111000010000111001001010111101000101100"; --    +422023   +2456108
      WHEN 1232 => Ti := "000100101110001100111000001011011000000110010000"; --   +1237816   +2982288
      WHEN 1233 => Ti := "001100011000010110001001111011001010110011011001"; --   +3245449   -1266471
      WHEN 1234 => Ti := "001011000101011100000100111110001100111010111011"; --   +2905860    -471365
      WHEN 1235 => Ti := "111111100101010100100100000010110011001001011100"; --    -109276    +733788
      WHEN 1236 => Ti := "000101100100000000011001110111100011101110110110"; --   +1458201   -2212938
      WHEN 1237 => Ti := "111011010010101111110001110100100100100100001000"; --   -1233935   -2995960
      WHEN 1238 => Ti := "111000101000100001111110000000001100001000011101"; --   -1931138     +49693
      WHEN 1239 => Ti := "110111000010101010111110110011101101101010001101"; --   -2348354   -3220851
      WHEN 1240 => Ti := "111010101101101100010110000001000011111000110010"; --   -1385706    +278066
      WHEN 1241 => Ti := "000000111111010001111000001001000010111011110001"; --    +259192   +2371313
      WHEN 1242 => Ti := "110011000010101111111000111100010000110000100110"; --   -3396616    -979930
      WHEN 1243 => Ti := "111010010100111111011001110110010011010001100100"; --   -1486887   -2542492
      WHEN 1244 => Ti := "110011000010000011000100000001010111001100000110"; --   -3399484    +357126
      WHEN 1245 => Ti := "110100111101111010001100000110111010111010111110"; --   -2892148   +1814206
      WHEN 1246 => Ti := "000111101001011101111110001010110011110010110101"; --   +2004862   +2833589
      WHEN 1247 => Ti := "111100110101010011100010111000101010011000110111"; --    -830238   -1923529
      WHEN 1248 => Ti := "000110110110100111010001111110110010001110010110"; --   +1796561    -318570
      WHEN 1249 => Ti := "001010011100001011110100001001101100100010011011"; --   +2736884   +2541723
      WHEN 1250 => Ti := "000011100000010010110100000001000110111111001101"; --    +918708    +290765
      WHEN 1251 => Ti := "000010101100111111010100111001101101101111101001"; --    +708564   -1647639
      WHEN 1252 => Ti := "000101010010010110101100000011110010101101000000"; --   +1385900    +994112
      WHEN 1253 => Ti := "000001100111001000100001001011101110111111111111"; --    +422433   +3076095
      WHEN 1254 => Ti := "111011111001110110011001110111000010001000001111"; --   -1073767   -2350577
      WHEN 1255 => Ti := "000110111011111101101101001001010010111000101011"; --   +1818477   +2436651
      WHEN 1256 => Ti := "001011000111111111010001000110010010010100010110"; --   +2916305   +1647894
      WHEN 1257 => Ti := "110101110011000000111010000111111101101011010111"; --   -2674630   +2087639
      WHEN 1258 => Ti := "110011101010010110100000110110010101111110011001"; --   -3234400   -2531431
      WHEN 1259 => Ti := "111110010010001101101011001011011100101111111000"; --    -449685   +3001336
      WHEN 1260 => Ti := "000011010101010010110000111000100000101100000000"; --    +873648   -1963264
      WHEN 1261 => Ti := "111011100000111100101001111000011000010010010110"; --   -1175767   -1997674
      WHEN 1262 => Ti := "000011101000000110000100000110110010101110001000"; --    +950660   +1780616
      WHEN 1263 => Ti := "110110111101000001010101001011101111011111111111"; --   -2371499   +3078143
      WHEN 1264 => Ti := "110111100011110100110001000011100011010110100001"; --   -2212559    +931233
      WHEN 1265 => Ti := "110100111110110000100110111110001001001010111010"; --   -2888666    -486726
      WHEN 1266 => Ti := "000110010111100000101100111101011010110001000010"; --   +1669164    -676798
      WHEN 1267 => Ti := "001000010011011011000001000110111101001010111111"; --   +2176705   +1823423
      WHEN 1268 => Ti := "111101011011100110111101000101000010001101011110"; --    -673347   +1319774
      WHEN 1269 => Ti := "000011011010111001001100000000000101001000011011"; --    +896588     +21019
      WHEN 1270 => Ti := "111010010010010010100101110101011101001110000011"; --   -1497947   -2763901
      WHEN 1271 => Ti := "111000111100010010000101110111111111000101011010"; --   -1850235   -2100902
      WHEN 1272 => Ti := "110011110110010011011000000011001110001111111111"; --   -3185448    +844799
      WHEN 1273 => Ti := "111011100011100011000100001100011000100000001110"; --   -1165116   +3246094
      WHEN 1274 => Ti := "000000100000111011010011001100011011110000001111"; --    +134867   +3259407
      WHEN 1275 => Ti := "000001101000101110111011110100101111100111011001"; --    +428987   -2950695
      WHEN 1276 => Ti := "110110101100010111101001111101111011000100011011"; --   -2439703    -544485
      WHEN 1277 => Ti := "110110111010101010111011111101100000010001000100"; --   -2381125    -654268
      WHEN 1278 => Ti := "111000100110111000010111111011000011101001110000"; --   -1937897   -1295760
      WHEN 1279 => Ti := "111001110011011000110011110100101010001101110000"; --   -1624525   -2972816
      WHEN 1280 => Ti := "001000111011001110011101000010100101011001010111"; --   +2339741    +677463
      WHEN 1281 => Ti := "000001111011111111000010111011110111101101010000"; --    +507842   -1082544
      WHEN 1282 => Ti := "000101110110100110111001001010111100000010111000"; --   +1534393   +2867384
      WHEN 1283 => Ti := "000111001101110001000001110011111110010011111001"; --   +1891393   -3152647
      WHEN 1284 => Ti := "110101000101000000101000000011100101111001101111"; --   -2863064    +941679
      WHEN 1285 => Ti := "000000011100110001101011110101111110000100101001"; --    +117867   -2629335
      WHEN 1286 => Ti := "111110001010011010011100000010101010101100100101"; --    -481636    +699173
      WHEN 1287 => Ti := "000100000101111100101001110011110110000111000011"; --   +1072937   -3186237
      WHEN 1288 => Ti := "111101110001011101011111001100011000000110101000"; --    -583841   +3244456
      WHEN 1289 => Ti := "111011110010101100110000110101010000010111100101"; --   -1103056   -2816539
      WHEN 1290 => Ti := "110101110001110111010011001000010101010101000111"; --   -2679341   +2184519
      WHEN 1291 => Ti := "000010000000111111000100001010011100111001000110"; --    +528324   +2739782
      WHEN 1292 => Ti := "110111110011000001101010000101100000010100000011"; --   -2150294   +1443075
      WHEN 1293 => Ti := "110100000110110011011110000011000011001001100010"; --   -3117858    +799330
      WHEN 1294 => Ti := "000001010111111011101000111010011010010011000111"; --    +360168   -1465145
      WHEN 1295 => Ti := "000011001101101001000111000011000100111001100010"; --    +842311    +806498
      WHEN 1296 => Ti := "000001000001110001111001001000110010011000011110"; --    +269433   +2303518
      WHEN 1297 => Ti := "000001101000111000100001000011110101010110101000"; --    +429601   +1004968
      WHEN 1298 => Ti := "111011010101111100100101001011110111110011001111"; --   -1220827   +3112143
      WHEN 1299 => Ti := "000011110111100110001010110100101000001101101111"; --   +1014154   -2981009
      WHEN 1300 => Ti := "000111010011111010101001111000100100100101101000"; --   +1916585   -1947288
      WHEN 1301 => Ti := "111001001110110101011001001000111101011110111100"; --   -1774247   +2348988
      WHEN 1302 => Ti := "111111100000111010111100001001110111100101101100"; --    -127300   +2586988
      WHEN 1303 => Ti := "000110100111100111001100000001101110110101110101"; --   +1735116    +454005
      WHEN 1304 => Ti := "000101110001101010000100110011110110100011110110"; --   +1514116   -3184394
      WHEN 1305 => Ti := "111010011100001001000011111111001001010001101100"; --   -1457597    -224148
      WHEN 1306 => Ti := "000011101001000010111000111110010000000100100011"; --    +954552    -458461
      WHEN 1307 => Ti := "001010101001110101100000110101100111100100100001"; --   +2792800   -2721503
      WHEN 1308 => Ti := "111000100001101011100001110011111101011010010011"; --   -1959199   -3156333
      WHEN 1309 => Ti := "000000110100001110100111000110100100100111101001"; --    +213927   +1722857
      WHEN 1310 => Ti := "110011000110101100101100111011101010010000011000"; --   -3380436   -1137640
      WHEN 1311 => Ti := "000101000000111001110010001010101001010101111110"; --   +1314418   +2790782
      WHEN 1312 => Ti := "000110110000000100000010111010010000111100101010"; --   +1769730   -1503446
      WHEN 1313 => Ti := "111000011010100001111000110100100101100000111011"; --   -1988488   -2992069
      WHEN 1314 => Ti := "000001000001010001111001111001100111111111100111"; --    +267385   -1671193
      WHEN 1315 => Ti := "110110101100100001001111110011111110011010010011"; --   -2439089   -3152237
      WHEN 1316 => Ti := "111100110011100110101110000001000101001011111111"; --    -837202    +283391
      WHEN 1317 => Ti := "001000101100110100110001111111000000010001101000"; --   +2280753    -261016
      WHEN 1318 => Ti := "111101100001011010001100110011110111010111000100"; --    -649588   -3181116
      WHEN 1319 => Ti := "000101111100111010001001110111010011000001111100"; --   +1560201   -2281348
      WHEN 1320 => Ti := "111100101111001101000110111100100011110111000111"; --    -855226    -901689
      WHEN 1321 => Ti := "111100001110101100111010110111011001101110110010"; --    -988358   -2253902
      WHEN 1322 => Ti := "111011000100111111101011111111111111101000011001"; --   -1290261      -1511
      WHEN 1323 => Ti := "000001001011011110110000111100111010000111001111"; --    +309168    -810545
      WHEN 1324 => Ti := "111110110000101101110111000101001100101101100010"; --    -324745   +1362786
      WHEN 1325 => Ti := "111000010111111000010001111100110100111010011010"; --   -1999343    -831846
      WHEN 1326 => Ti := "110110111110111110001001001100110011111101001100"; --   -2363511   +3358540
      WHEN 1327 => Ti := "111110101000101101110100111100100111110111001001"; --    -357516    -885303
      WHEN 1328 => Ti := "001000001011000111110001111000101110100010011110"; --   +2142705   -1906530
      WHEN 1329 => Ti := "000101000000000011011000001010010010011111011100"; --   +1310936   +2697180
      WHEN 1330 => Ti := "000101000100000110100111111110011010000100100111"; --   +1327527    -417497
      WHEN 1331 => Ti := "111111010101000100011110111010101011000000000000"; --    -175842   -1396736
      WHEN 1332 => Ti := "111111000011001010110001110111110100101110111100"; --    -249167   -2143300
      WHEN 1333 => Ti := "111101110010000000101100111011101010010000011000"; --    -581588   -1137640
      WHEN 1334 => Ti := "111110100100010100001100110011110111100011110111"; --    -375540   -3180297
      WHEN 1335 => Ti := "111011100001010110010000111011000000000110100010"; --   -1174128   -1310302
      WHEN 1336 => Ti := "000001001001000101001001110011110011011010001111"; --    +299337   -3197297
      WHEN 1337 => Ti := "000110101100010111001110001000111111001011110000"; --   +1754574   +2355952
      WHEN 1338 => Ti := "000001000100101110101101000011010111100011010000"; --    +281517    +882896
      WHEN 1339 => Ti := "001100000001110010110100000100100100110000100000"; --   +3153076   +1199136
      WHEN 1340 => Ti := "001010110010000101100011111111100001011110101000"; --   +2826595    -125016
      WHEN 1341 => Ti := "000011101101101001010011000100111110010011110110"; --    +973395   +1303798
      WHEN 1342 => Ti := "001010001100010101010101000110010001001010101111"; --   +2671957   +1643183
      WHEN 1343 => Ti := "111101000111001010000011000001011101110101101111"; --    -757117    +384367
      WHEN 1344 => Ti := "000111011000010001000100111101000101000100000111"; --   +1934404    -765689
      WHEN 1345 => Ti := "111010000111111000111011111000010010101011111010"; --   -1540549   -2020614
      WHEN 1346 => Ti := "111100110110110011100011110101001110010001001010"; --    -824093   -2825142
      WHEN 1347 => Ti := "111110001100101101101001111011110001010110110100"; --    -472215   -1108556
      WHEN 1348 => Ti := "111110101110000001000011110101000110110111100001"; --    -335805   -2855455
      WHEN 1349 => Ti := "110101000000100011110100000000000101011000011011"; --   -2881292     +22043
      WHEN 1350 => Ti := "110110101000010111100111000111011110110111111111"; --   -2456089   +1961471
      WHEN 1351 => Ti := "000111111101100100011111000100000110010110101110"; --   +2087199   +1074606
      WHEN 1352 => Ti := "111000101010101110110010111110000101110001010010"; --   -1922126    -500654
      WHEN 1353 => Ti := "000110100011110111001010001001010000001011110110"; --   +1719754   +2425590
      WHEN 1354 => Ti := "110101000000011101011010111011110001110000011011"; --   -2881702   -1106917
      WHEN 1355 => Ti := "111000110100110101001111110100110111110001000010"; --   -1880753   -2917310
      WHEN 1356 => Ti := "111101101010111010010000000000011100010101010110"; --    -610672    +116054
      WHEN 1357 => Ti := "111111110000110111110101000010001010100010110011"; --     -61963    +567475
      WHEN 1358 => Ti := "111101111010000111001001001010110101101100011100"; --    -548407   +2841372
      WHEN 1359 => Ti := "000001011110010010000100111000110101001100000111"; --    +386180   -1879289
      WHEN 1360 => Ti := "000000110110001110101000001010101000001001001011"; --    +222120   +2785867
      WHEN 1361 => Ti := "111000000111011011011000000010110000011111110100"; --   -2066728    +722932
      WHEN 1362 => Ti := "111110100101000000111111000011011110110000000110"; --    -372673    +912390
      WHEN 1363 => Ti := "111010111011111001001110000111111011101110100100"; --   -1327538   +2079652
      WHEN 1364 => Ti := "000000011111110100111001000010000010100010110000"; --    +130361    +534704
      WHEN 1365 => Ti := "001011101101111001000110000100101000100000100001"; --   +3071558   +1214497
      WHEN 1366 => Ti := "111010011111101100010001110110101101100001101110"; --   -1443055   -2434962
      WHEN 1367 => Ti := "110011000110011001011111110100001111101101100110"; --   -3381665   -3081370
      WHEN 1368 => Ti := "110110100110010100011010111101100001100100010001"; --   -2464486    -648943
      WHEN 1369 => Ti := "000010111101100101110100110111111101000101011001"; --    +776564   -2109095
      WHEN 1370 => Ti := "001010010000111011110000110011110101001010010000"; --   +2690800   -3190128
      WHEN 1371 => Ti := "001001001101011011010111000110110111000100100011"; --   +2414295   +1798435
      WHEN 1372 => Ti := "111111101101010111110100111100101010010111001010"; --     -76300    -875062
      WHEN 1373 => Ti := "111101011101010011110001000001111101010101111011"; --    -666383    +513403
      WHEN 1374 => Ti := "110111010100000111111000000111101110101011010010"; --   -2276872   +2026194
      WHEN 1375 => Ti := "000000110000000001110010111001100100101111100110"; --    +196722   -1684506
      WHEN 1376 => Ti := "000101000011111001110011111011110111111101010000"; --   +1326707   -1081520
      WHEN 1377 => Ti := "000110100000110000110000111110101000110111111001"; --   +1707056    -356871
      WHEN 1378 => Ti := "110100011010010000011000111111011000011110100100"; --   -3038184    -161884
      WHEN 1379 => Ti := "001010110001011111001001000000100111000101011010"; --   +2824137    +160090
      WHEN 1380 => Ti := "000011011101110110000000111110111011001011001101"; --    +908672    -281907
      WHEN 1381 => Ti := "111001101000011000101111111000110111000010100010"; --   -1669585   -1871710
      WHEN 1382 => Ti := "001100100010101100100111000111001010100100101011"; --   +3287847   +1878315
      WHEN 1383 => Ti := "111000110001011011100111111101111001100100011010"; --   -1894681    -550630
      WHEN 1384 => Ti := "001000100111011011001001111000001101101011111001"; --   +2258633   -2041095
      WHEN 1385 => Ti := "000011110101001111101111111111010000001011010100"; --   +1004527    -195884
      WHEN 1386 => Ti := "111011011010110110001101110011101110111101011010"; --   -1200755   -3215526
      WHEN 1387 => Ti := "001100011010000010111101110111100101110101010000"; --   +3252413   -2204336
      WHEN 1388 => Ti := "000000011000001011010000001100111000111101001110"; --     +99024   +3379022
      WHEN 1389 => Ti := "110100111011010011110010001001000111000101011001"; --   -2902798   +2388313
      WHEN 1390 => Ti := "001001001100011110100011000001010110000101101100"; --   +2410403    +352620
      WHEN 1391 => Ti := "111101100100110000100111000100111100111101011100"; --    -635865   +1298268
      WHEN 1392 => Ti := "000101010011001101000110000010100010000010111100"; --   +1389382    +663740
      WHEN 1393 => Ti := "111010011100000010101001000100111001001010001110"; --   -1458007   +1282702
      WHEN 1394 => Ti := "000010111011111111011010001001100010011111001010"; --    +770010   +2500554
      WHEN 1395 => Ti := "000011101111010010111010111110011101100001011011"; --    +980154    -403365
      WHEN 1396 => Ti := "000001000110101110101110001001101010110101100111"; --    +289710   +2534759
      WHEN 1397 => Ti := "110111010010010100101010110110101110011000001000"; --   -2284246   -2431480
      WHEN 1398 => Ti := "000011001001100010101100111100000010111101010100"; --    +825516   -1036460
      WHEN 1399 => Ti := "111100000000100000000010001010101101110110000000"; --   -1046526   +2809216
      WHEN 1400 => Ti := "000011100110010010110111111110101010100100101101"; --    +943287    -349907
      WHEN 1401 => Ti := "111000010011000101000010110011101100110011110011"; --   -2019006   -3224333
      WHEN 1402 => Ti := "001010010000101011110000000001010010110010011110"; --   +2689776    +339102
      WHEN 1403 => Ti := "111000110110010010000011001000001000000101000010"; --   -1874813   +2130242
      WHEN 1404 => Ti := "000011001010001001000110000111011011011011001011"; --    +827974   +1947339
      WHEN 1405 => Ti := "111000101100111011100110111001111110011111110000"; --   -1913114   -1579024
      WHEN 1406 => Ti := "000000101110011110100101111001101100011001001111"; --    +190373   -1653169
      WHEN 1407 => Ti := "001000001011011010111110000110100111101110000100"; --   +2143934   +1735556
      WHEN 1408 => Ti := "000110110110001010011110110100010011010100000001"; --   +1794718   -3066623
      WHEN 1409 => Ti := "110110101000001110000001001100000100110110100000"; --   -2456703   +3165600
      WHEN 1410 => Ti := "001001001000101110100010110011010110011101010001"; --   +2395042   -3315887
      WHEN 1411 => Ti := "111100101010100110101011000100100010101101010010"; --    -874069   +1190738
      WHEN 1412 => Ti := "000110111001011101101100111101110001110100011000"; --   +1808236    -582376
      WHEN 1413 => Ti := "001010110100001011111101110101110010000100100101"; --   +2835197   -2678491
      WHEN 1414 => Ti := "001000101100110111111110111100100100000011111010"; --   +2280958    -900870
      WHEN 1415 => Ti := "000111000010011010100011001000010110011011100001"; --   +1844899   +2189025
      WHEN 1416 => Ti := "000011101000001100011110111000100101010010011011"; --    +951070   -1944421
      WHEN 1417 => Ti := "000011011111101111100111000111011101010001100101"; --    +916455   +1954917
      WHEN 1418 => Ti := "111111110000110100101001000110010100001010110000"; --     -62167   +1655472
      WHEN 1419 => Ti := "000101110001001101010001111101100001000100010001"; --   +1512273    -650991
      WHEN 1420 => Ti := "000101111011101010001000000000001011111000011101"; --   +1555080     +48669
      WHEN 1421 => Ti := "000010100000111100000011111010111010100000000110"; --    +659203   -1333242
      WHEN 1422 => Ti := "111111000101111101111111001001111110110101101110"; --    -237697   +2616686
      WHEN 1423 => Ti := "001011001100001111010011000111110101011110100001"; --   +2933715   +2054049
      WHEN 1424 => Ti := "001001011000011000001110111110000110000100011111"; --   +2459150    -499425
      WHEN 1425 => Ti := "000101000001000000001100000001111100010010101110"; --   +1314828    +509102
      WHEN 1426 => Ti := "000110110010100100000011001011110101010011001110"; --   +1779971   +3101902
      WHEN 1427 => Ti := "000000011000101011010000000000010011101110111010"; --    +101072     +80826
      WHEN 1428 => Ti := "000011000111110101111000110100010111000100000011"; --    +818552   -3051261
      WHEN 1429 => Ti := "000111111100011110000101111110011000111110001101"; --   +2082693    -422003
      WHEN 1430 => Ti := "000001111110100010010000111010010100100110010010"; --    +518288   -1488494
      WHEN 1431 => Ti := "111110011111011101110000000010000011101111100100"; --    -395408    +539620
      WHEN 1432 => Ti := "000101100101100110110011001011010001101100100111"; --   +1464755   +2956071
      WHEN 1433 => Ti := "111100100011011001110101111101011110011010101010"; --    -903563    -661846
      WHEN 1434 => Ti := "111000111010010101010001000011110011011101000001"; --   -1858223    +997185
      WHEN 1435 => Ti := "110111111111101110100010000111001110010001011111"; --   -2098270   +1893471
      WHEN 1436 => Ti := "000000111110101011011110111011110111100011101010"; --    +256734   -1083158
      WHEN 1437 => Ti := "110011010010110011001010110110010001110100110001"; --   -3330870   -2548431
      WHEN 1438 => Ti := "111001011110011000101011111100001101101010001100"; --   -1710549    -992628
      WHEN 1439 => Ti := "111110110110000001000110111100010000000111000000"; --    -303034    -982592
      WHEN 1440 => Ti := "000110111111000000111011001010011010100010101100"; --   +1830971   +2730156
      WHEN 1441 => Ti := "111101001000000110110110111110101001100111111001"; --    -753226    -353799
      WHEN 1442 => Ti := "000010111000001111011001000101111110110111011011"; --    +754649   +1568219
      WHEN 1443 => Ti := "110100001000010000010010111100110100010000110100"; --   -3111918    -834508
      WHEN 1444 => Ti := "111000000011111110100011110111010100100001111101"; --   -2080861   -2275203
      WHEN 1445 => Ti := "110110011010000100010101110110100000000100110110"; --   -2514667   -2490058
      WHEN 1446 => Ti := "110100100011110011101001111110001000010001010011"; --   -2999063    -490413
      WHEN 1447 => Ti := "000111110011011010110101000111000110010111110110"; --   +2045621   +1861110
      WHEN 1448 => Ti := "000000110000011000001100000000000011000010000000"; --    +198156     +12416
      WHEN 1449 => Ti := "001000001101000001011000110110010011111110011000"; --   +2150488   -2539624
      WHEN 1450 => Ti := "000000010010011000000001111000010111011011111100"; --     +75265   -2001156
      WHEN 1451 => Ti := "001000010111010111110110001011111001100011001111"; --   +2192886   +3119311
      WHEN 1452 => Ti := "000000100101010001101110001001100101011000110010"; --    +152686   +2512434
      WHEN 1453 => Ti := "111001100100110010010100000000110100111111000110"; --   -1684332    +217030
      WHEN 1454 => Ti := "000101110110101101010011111110011001010111110011"; --   +1534803    -420365
      WHEN 1455 => Ti := "000010100100100010011110110101001000001101111011"; --    +673950   -2849925
      WHEN 1456 => Ti := "110100001000110011011111110100100100000111010100"; --   -3109665   -2997804
      WHEN 1457 => Ti := "000100000110001100101001110111111101001011110010"; --   +1073961   -2108686
      WHEN 1458 => Ti := "001011100101100010101001111000110011110010100000"; --   +3037353   -1885024
      WHEN 1459 => Ti := "111101111011011101100011001001000111111011110011"; --    -542877   +2391795
      WHEN 1460 => Ti := "111011111111111100110101000001010111011111010011"; --   -1048779    +358355
      WHEN 1461 => Ti := "111000010101100101000011001000000100111011011010"; --   -2008765   +2117338
      WHEN 1462 => Ti := "000110110101001101101011110100110010100001000000"; --   +1790827   -2938816
      WHEN 1463 => Ti := "001001001100111110100011110111100001101000011011"; --   +2412451   -2221541
      WHEN 1464 => Ti := "000000011010101011010001110111011001111000011000"; --    +109265   -2253288
      WHEN 1465 => Ti := "111111001011001010110100001001101110100010011011"; --    -216396   +2549915
      WHEN 1466 => Ti := "110100011110000011100111111001110011111001010010"; --   -3022617   -1622446
      WHEN 1467 => Ti := "111101010011010110111010110110001100101110010101"; --    -707142   -2569323
      WHEN 1468 => Ti := "001011011011001000111111110110000010001110010001"; --   +2994751   -2612335
      WHEN 1469 => Ti := "110111111000101011010010001100111010101101001110"; --   -2127150   +3386190
      WHEN 1470 => Ti := "110100100111000110110111001000111100000010001000"; --   -2985545   +2343048
      WHEN 1471 => Ti := "110110100110010111100110000111101110001110011110"; --   -2464282   +2024350
      WHEN 1472 => Ti := "001100100001101111110011001000101010000010000010"; --   +3283955   +2269314
      WHEN 1473 => Ti := "110011000011011001011110110100011010100111010001"; --   -3393954   -3036719
      WHEN 1474 => Ti := "000011000101110101110111111000111010111100001010"; --    +810359   -1855734
      WHEN 1475 => Ti := "000100100111010110011100000101000101011101011111"; --   +1209756   +1333087
      WHEN 1476 => Ti := "000110000000110110111101111110000000001010110111"; --   +1576381    -523593
      WHEN 1477 => Ti := "111101011101101010001011000111011101111110011000"; --    -664949   +1957784
      WHEN 1478 => Ti := "111111111110000111111010111011111010010011101011"; --      -7686   -1071893
      WHEN 1479 => Ti := "110110100001001101111110000100001100101001111101"; --   -2485378   +1100413
      WHEN 1480 => Ti := "001010010000000101010110000010101001111111110010"; --   +2687318    +696306
      WHEN 1481 => Ti := "000111110011010111101000111001110111110010111010"; --   +2045416   -1606470
      WHEN 1482 => Ti := "001000000010110100100001000001111100010101111010"; --   +2108705    +509306
      WHEN 1483 => Ti := "110111101001000111111111000001100101011000111111"; --   -2190849    +415295
      WHEN 1484 => Ti := "001000111110110100111000111110101110110111111011"; --   +2354488    -332293
      WHEN 1485 => Ti := "000100110000101001101100000100000110011001111011"; --   +1247852   +1074811
      WHEN 1486 => Ti := "000011101110101001010011111000001111011000101100"; --    +977491   -2034132
      WHEN 1487 => Ti := "111011111101101100110100000000011111000101010111"; --   -1057996    +127319
      WHEN 1488 => Ti := "000110001110100000101001000011100101111100111100"; --   +1632297    +941884
      WHEN 1489 => Ti := "001010010101010101011000001011011000110011000011"; --   +2708824   +2985155
      WHEN 1490 => Ti := "000101111110011101010110111110111011001000000000"; --   +1566550    -282112
      WHEN 1491 => Ti := "111100100111100000010000000111110000011110011111"; --    -886768   +2033567
      WHEN 1492 => Ti := "000111100101100001001001111100101111000111001011"; --   +1988681    -855605
      WHEN 1493 => Ti := "110110010100001101111001110011011011101010000110"; --   -2538631   -3294586
      WHEN 1494 => Ti := "111011001010001100100001111011011111111101000111"; --   -1268959   -1179833
      WHEN 1495 => Ti := "000100011000111001100011111011100100010110101111"; --   +1150563   -1161809
      WHEN 1496 => Ti := "000100101111010000000101001010010011100010101001"; --   +1242117   +2701481
      WHEN 1497 => Ti := "111100011010011100111111000000000110101110110101"; --    -940225     +27573
      WHEN 1498 => Ti := "110100110010010000100001001000001010101110101001"; --   -2939871   +2141097
      WHEN 1499 => Ti := "001100001101111100011111000111000110111011000011"; --   +3202847   +1863363
      WHEN 1500 => Ti := "110100101111001010000111000101001011011101100010"; --   -2952569   +1357666
      WHEN 1501 => Ti := "000100010100111100101111111010010101011111111000"; --   +1134383   -1484808
      WHEN 1502 => Ti := "111000011000101011011110001100101101110011100011"; --   -1996066   +3333347
      WHEN 1503 => Ti := "110100011111100110110100111100101011010111001010"; --   -3016268    -870966
      WHEN 1504 => Ti := "111000000111101011011000111001011110101111100100"; --   -2065704   -1709084
      WHEN 1505 => Ti := "001011000100000010011101111110100111110111111001"; --   +2900125    -360967
      WHEN 1506 => Ti := "000100110100100110100001000001000001011011111110"; --   +1264033    +268030
      WHEN 1507 => Ti := "000001100100011110111001111000111111101100001011"; --    +411577   -1836277
      WHEN 1508 => Ti := "000110001100101101011011111101110111110111100111"; --   +1624923    -557593
      WHEN 1509 => Ti := "000111011011100100010011110101001000001101111011"; --   +1947923   -2849925
      WHEN 1510 => Ti := "000001001011100101001010001100010111001001110100"; --    +309578   +3240564
      WHEN 1511 => Ti := "110101000010011010001110111100111001010100000010"; --   -2873714    -813822
      WHEN 1512 => Ti := "000011111101011111110011000001010000100101101010"; --   +1038323    +330090
      WHEN 1513 => Ti := "000100111100011001110000000000001011101110110111"; --   +1295984     +48055
      WHEN 1514 => Ti := "111011101011011111111010000001011111011100001001"; --   -1132550    +390921
      WHEN 1515 => Ti := "110111000011011110001011111101011011010001000010"; --   -2345077    -674750
      WHEN 1516 => Ti := "110111110001101000000011110101010001111101111111"; --   -2156029   -2809985
      WHEN 1517 => Ti := "110101000111100000101001111010110001111100110110"; --   -2852823   -1368266
      WHEN 1518 => Ti := "000101010111011101000111000100010111010011101000"; --   +1406791   +1144040
      WHEN 1519 => Ti := "000010110100101100001010000011111101000011011110"; --    +740106   +1036510
      WHEN 1520 => Ti := "110011011111011001101001001000110100111110111001"; --   -3279255   +2314169
      WHEN 1521 => Ti := "000011111110010110001100000111000101010001011100"; --   +1041804   +1856604
      WHEN 1522 => Ti := "110111011010001011000111001100100111111101000111"; --   -2252089   +3309383
      WHEN 1523 => Ti := "001001100000001011011110110111110110110101010110"; --   +2491102   -2134698
      WHEN 1524 => Ti := "000001101110110101010111001100000111101100111011"; --    +453975   +3177275
      WHEN 1525 => Ti := "001001010101010101000000111001101101011111101001"; --   +2446656   -1648663
      WHEN 1526 => Ti := "001000011010100001011101111000000110011000101001"; --   +2205789   -2070999
      WHEN 1527 => Ti := "111110101100111010101001111000001110111111000110"; --    -340311   -2035770
      WHEN 1528 => Ti := "111100110011001001111011111110011011000111110100"; --    -839045    -413196
      WHEN 1529 => Ti := "111101010100100000100001001000010000110101000101"; --    -702431   +2166085
      WHEN 1530 => Ti := "111110100000011101110001111010000111101001011001"; --    -391311   -1541543
      WHEN 1531 => Ti := "000001110010011110111110111000110010111100000111"; --    +468926   -1888505
      WHEN 1532 => Ti := "000010011000000010011001111000100011000010011010"; --    +622745   -1953638
      WHEN 1533 => Ti := "001001101010101000010101000111110010101000000111"; --   +2533909   +2042375
      WHEN 1534 => Ti := "111110001111110111010001000001001100100010011100"; --    -459311    +313500
      WHEN 1535 => Ti := "001010011000010101011001001000010111110001111011"; --   +2721113   +2194555
      WHEN 1536 => Ti := "000100000001001111110100110100001000110000110000"; --   +1053684   -3109840
      WHEN 1537 => Ti := "000100100110011001101000001000000111101011011011"; --   +1205864   +2128603
      WHEN 1538 => Ti := "110110010100100001000110111001100010000101111111"; --   -2537402   -1695361
      WHEN 1539 => Ti := "111110011100011101101111110100001100101101100101"; --    -407697   -3093659
      WHEN 1540 => Ti := "110100011101110110110011001001011000011111000110"; --   -3023437   +2459590
      WHEN 1541 => Ti := "001000100011101110010100111111001000110001101011"; --   +2243476    -226197
      WHEN 1542 => Ti := "110100110101110000100011000101111011010100001101"; --   -2925533   +1553677
      WHEN 1543 => Ti := "111110110011110100010010111011001111100000001110"; --    -312046   -1247218
      WHEN 1544 => Ti := "111000001000101011011000001001100000011111001001"; --   -2061608   +2492361
      WHEN 1545 => Ti := "110101011110011101100101000100000110010000010100"; --   -2758811   +1074196
      WHEN 1546 => Ti := "111111110110010100101011111011110111001010000011"; --     -39637   -1084797
      WHEN 1547 => Ti := "000011101001100110000101110111110111111011110000"; --    +956805   -2130192
      WHEN 1548 => Ti := "111111001101111110000010110110000101001110010010"; --    -204926   -2600046
      WHEN 1549 => Ti := "110101010011000111000111000001010100100010011111"; --   -2805305    +346271
      WHEN 1550 => Ti := "001010100111011011111000001001001101111011110110"; --   +2782968   +2416374
      WHEN 1551 => Ti := "111100001100100000000110111111111110111110110011"; --    -997370      -4173
      WHEN 1552 => Ti := "111100100101011101000011001000010100011110101101"; --    -895165   +2181037
      WHEN 1553 => Ti := "000011101010111001010010110101111001000001011010"; --    +962130   -2650022
      WHEN 1554 => Ti := "000111101111010001001101000011100011101100111011"; --   +2028621    +932667
      WHEN 1555 => Ti := "001011001110111000111010111011011110100011100000"; --   +2944570   -1185568
      WHEN 1556 => Ti := "000110010010011010010001111011100100001001111100"; --   +1648273   -1162628
      WHEN 1557 => Ti := "111000110101011000011100111010100011111001100100"; --   -1878500   -1425820
      WHEN 1558 => Ti := "111110011100010111010110111010101001001001100110"; --    -408106   -1404314
      WHEN 1559 => Ti := "111001111111011111010001111101111110011010110110"; --   -1574959    -530762
      WHEN 1560 => Ti := "111001010000000101011001000001011010011100000111"; --   -1769127    +370439
      WHEN 1561 => Ti := "111110001001001101101000001001110110001100000101"; --    -486552   +2581253
      WHEN 1562 => Ti := "001001011111001000010001110100100001010100000110"; --   +2486801   -3009274
      WHEN 1563 => Ti := "111011000100011001010010111101010100001101110011"; --   -1292718    -703629
      WHEN 1564 => Ti := "000110100101011101100101111000111111011111011000"; --   +1726309   -1837096
      WHEN 1565 => Ti := "000101110000001101010001001011010101000011000010"; --   +1508177   +2969794
      WHEN 1566 => Ti := "001100011100101111110001000110011011101010110011"; --   +3263473   +1686195
      WHEN 1567 => Ti := "001010000110101011101100111110011100110100101000"; --   +2648812    -406232
      WHEN 1568 => Ti := "110111010001010001011101000011000100111100101111"; --   -2288547    +806703
      WHEN 1569 => Ti := "111000101101110101001100001000100011100101001100"; --   -1909428   +2242892
      WHEN 1570 => Ti := "000101110101110011101100111101101101000100010110"; --   +1531116    -601834
      WHEN 1571 => Ti := "000001111001000010001110000101100011000100000100"; --    +495758   +1454340
      WHEN 1572 => Ti := "110011000100011111111000001100100101000011100000"; --   -3389448   +3297504
      WHEN 1573 => Ti := "000001111001010101011011001011100010101100101101"; --    +496987   +3025709
      WHEN 1574 => Ti := "111110000000000111001011111111000011101110011101"; --    -523829    -246883
      WHEN 1575 => Ti := "000010011110111000110110111100011111010011111001"; --    +650806    -920327
      WHEN 1576 => Ti := "111101110100111101100001000010101001100110001011"; --    -569503    +694667
      WHEN 1577 => Ti := "110101101001110000110110110011101010011010001011"; --   -2712522   -3234165
      WHEN 1578 => Ti := "111001001100101011110010000010101101001100100110"; --   -1783054    +709414
      WHEN 1579 => Ti := "110100000100111001110111110110001011010100101110"; --   -3125641   -2575058
      WHEN 1580 => Ti := "110111111101001110100001111101001011110100001001"; --   -2108511    -738039
      WHEN 1581 => Ti := "001001100011100101000101110100001010110000110001"; --   +2505029   -3101647
      WHEN 1582 => Ti := "000110100001110011111101111010000011000010111110"; --   +1711357   -1560386
      WHEN 1583 => Ti := "110011100010000011010000000001110100111001000100"; --   -3268400    +478788
      WHEN 1584 => Ti := "001000100011101110010100111001010100010101111001"; --   +2243476   -1751687
      WHEN 1585 => Ti := "110101101010110111010000001001000100010101011000"; --   -2708016   +2377048
      WHEN 1586 => Ti := "000101001101011101000100000101011000001101100110"; --   +1365828   +1409894
      WHEN 1587 => Ti := "110101010000010111000110110100101010100000111101"; --   -2816570   -2971587
      WHEN 1588 => Ti := "001010101101000010010100001010010100111001000011"; --   +2805908   +2707011
      WHEN 1589 => Ti := "111111011110001110001000111100000010000011101110"; --    -138360   -1040146
      WHEN 1590 => Ti := "000110101100101101100111000110011000001101111110"; --   +1756007   +1672062
      WHEN 1591 => Ti := "000100111010010000001001110110110101110001110001"; --   +1287177   -2401167
      WHEN 1592 => Ti := "111101111100011101100011000000111010111111001000"; --    -538781    +241608
      WHEN 1593 => Ti := "000111111011111010111000111001010011101001000110"; --   +2080440   -1754554
      WHEN 1594 => Ti := "000000110001010101000000110101110100011110001100"; --    +202048   -2668660
      WHEN 1595 => Ti := "001000010011101011000001000110101101110111101101"; --   +2177729   +1760749
      WHEN 1596 => Ti := "111010000001000010011111001000111101101110111100"; --   -1568609   +2350012
      WHEN 1597 => Ti := "000011001111010010101110000001011001100101101101"; --    +849070    +366957
      WHEN 1598 => Ti := "000010110101011111011000111100011110001010010010"; --    +743384    -925038
      WHEN 1599 => Ti := "000101100001000011100101001100001010110000001001"; --   +1446117   +3189769
      WHEN 1600 => Ti := "001100001000001001010000001010010110011001000100"; --   +3179088   +2713156
      WHEN 1601 => Ti := "110011101010011001101101000100011000011101001110"; --   -3234195   +1148750
      WHEN 1602 => Ti := "001000000001110111101110000010011000101100011111"; --   +2104814    +625439
      WHEN 1603 => Ti := "000101110000100011101010111011111000110011101010"; --   +1509610   -1078038
      WHEN 1604 => Ti := "111101110111000011111011000000010100000101010011"; --    -560901     +82259
      WHEN 1605 => Ti := "000001010010111000011001110011100101110000100011"; --    +339481   -3253213
      WHEN 1606 => Ti := "111111101101100111110100000001011010000010100001"; --     -75276    +368801
      WHEN 1607 => Ti := "111011100000011001011100001010101011111111100110"; --   -1178020   +2801638
      WHEN 1608 => Ti := "000101101011111010000010111010010101011111111000"; --   +1490562   -1484808
      WHEN 1609 => Ti := "111011010100100010111110111100111011101101101010"; --   -1226562    -803990
      WHEN 1610 => Ti := "001100011000011100100011000001010001011100000100"; --   +3245859    +333572
      WHEN 1611 => Ti := "111000100101101000010110001010011000110101111000"; --   -1943018   +2723192
      WHEN 1612 => Ti := "111010101001001100010100111001110101100010111001"; --   -1404140   -1615687
      WHEN 1613 => Ti := "110110001000100001000010001001011000001000101101"; --   -2586558   +2458157
      WHEN 1614 => Ti := "111000111100111011101100001010000111000010100101"; --   -1847572   +2650277
      WHEN 1615 => Ti := "000001000101011000010100001001111011100101101101"; --    +284180   +2603373
      WHEN 1616 => Ti := "001011010000100101101110111001011110010101111101"; --   +2951534   -1710723
      WHEN 1617 => Ti := "000110001110100000101001111110101010000001100000"; --   +1632297    -352160
      WHEN 1618 => Ti := "111110000100110111001101110011101110110111000000"; --    -504371   -3215936
      WHEN 1619 => Ti := "111011000001101100011101000101011110001010011100"; --   -1303779   +1434268
      WHEN 1620 => Ti := "110111101000000100110010000100011100110000011101"; --   -2195150   +1166365
      WHEN 1621 => Ti := "111110010010111101101100110111010111111011100100"; --    -446612   -2261276
      WHEN 1622 => Ti := "001010101000001111000110111000001001110010010001"; --   +2786246   -2057071
      WHEN 1623 => Ti := "000111101101000100011001001100111000011101001101"; --   +2019609   +3376973
      WHEN 1624 => Ti := "000001111011011111000010110111011001100101001011"; --    +505794   -2254517
      WHEN 1625 => Ti := "111101010110000000100010001011000110001111101111"; --    -696286   +2909167
      WHEN 1626 => Ti := "110101110011110111010100001001010001001011110111"; --   -2671148   +2429687
      WHEN 1627 => Ti := "111001110000001000110010111010001111101111110110"; --   -1637838   -1508362
      WHEN 1628 => Ti := "111011101110000110010100000100100000101101010010"; --   -1121900   +1182546
      WHEN 1629 => Ti := "111111111110010001100001001100110110110011100110"; --      -7071   +3370214
      WHEN 1630 => Ti := "000001010000101011100101000011010111011100110110"; --    +330469    +882486
      WHEN 1631 => Ti := "000001101010110010001000000101001010111101100001"; --    +437384   +1355617
      WHEN 1632 => Ti := "001001101000101011100001111010110011010011010000"; --   +2525921   -1362736
      WHEN 1633 => Ti := "110100111000111010001010001100110110010110110011"; --   -2912630   +3368371
      WHEN 1634 => Ti := "110111111011110001101101001001001110100101011100"; --   -2114451   +2419036
      WHEN 1635 => Ti := "110111000110000001011001111111101010111110101011"; --   -2334631     -86101
      WHEN 1636 => Ti := "000011111000100110001010000011110101100110101000"; --   +1018250   +1005992
      WHEN 1637 => Ti := "000111110011100111101000000011101111010000001100"; --   +2046440    +979980
      WHEN 1638 => Ti := "000011011011001001001100001001110100101100000100"; --    +897612   +2575108
      WHEN 1639 => Ti := "001011101110111100010011001001011110111000101111"; --   +3075859   +2485807
      WHEN 1640 => Ti := "110011100011101001101010001011000001001111101110"; --   -3261846   +2888686
      WHEN 1641 => Ti := "001001001000100001101111110100010110100111001111"; --   +2394223   -3053105
      WHEN 1642 => Ti := "000100011100011100110001001001001101101000101001"; --   +1165105   +2415145
      WHEN 1643 => Ti := "000001011011101011101001000110100011010111101001"; --    +375529   +1717737
      WHEN 1644 => Ti := "111001100001101111000110000001101100001111011011"; --   -1696826    +443355
      WHEN 1645 => Ti := "001100000101100110000010000011110010110000001101"; --   +3168642    +994317
      WHEN 1646 => Ti := "001000001001000001010111111001011100101100010110"; --   +2134103   -1717482
      WHEN 1647 => Ti := "111101000110010110110101001011111100100110011101"; --    -760395   +3131805
      WHEN 1648 => Ti := "000101010101100110101101000000000010011011100110"; --   +1399213      +9958
      WHEN 1649 => Ti := "000111111111001110000110000111111010011000001001"; --   +2093958   +2074121
      WHEN 1650 => Ti := "110011110010010000001001001001110111111111010010"; --   -3202039   +2588626
      WHEN 1651 => Ti := "110110011001000111100010110110010110000001100101"; --   -2518558   -2531227
      WHEN 1652 => Ti := "110101101101011101101011110101111111000001011101"; --   -2697365   -2625443
      WHEN 1653 => Ti := "111100110000011001111010001100001111010011011000"; --    -850310   +3208408
      WHEN 1654 => Ti := "000000011110111000000110000110011010111101111111"; --    +126470   +1683327
      WHEN 1655 => Ti := "110111011011000100101101110110111100011011011010"; --   -2248403   -2373926
      WHEN 1656 => Ti := "001001000011100001101101000101101100101101101110"; --   +2373741   +1493870
      WHEN 1657 => Ti := "000001000001010001111001000000011101101000100100"; --    +267385    +121380
      WHEN 1658 => Ti := "000110110111000000111000111010000111001001011001"; --   +1798200   -1543591
      WHEN 1659 => Ti := "111001010000011011110011111101001010000111010101"; --   -1767693    -745003
      WHEN 1660 => Ti := "000100010110001100101111000111101011110100110111"; --   +1139503   +2014519
      WHEN 1661 => Ti := "000110100110110011111111110110111100011000001101"; --   +1731839   -2374131
      WHEN 1662 => Ti := "000001001011000101001001111011001010011100111111"; --    +307529   -1267905
      WHEN 1663 => Ti := "110110110011110001010010111101000111000111010100"; --   -2409390    -757292
      WHEN 1664 => Ti := "110110110110000111101100000101010010011101100100"; --   -2399764   +1386340
      WHEN 1665 => Ti := "001000101001011110010110001100110011100011100101"; --   +2267030   +3356901
      WHEN 1666 => Ti := "110111000000100111110000000111000101000111110101"; --   -2356752   +1855989
      WHEN 1667 => Ti := "000010111100111111011010111001010110001111100001"; --    +774106   -1743903
      WHEN 1668 => Ti := "000000111111011110101011110110011001100001100111"; --    +260011   -2516889
      WHEN 1669 => Ti := "001001101011011011100010111011101000010110110001"; --   +2537186   -1145423
      WHEN 1670 => Ti := "000101110010010000011110001000010110101110101110"; --   +1516574   +2190254
      WHEN 1671 => Ti := "111011011010001100100111000010111011010110010010"; --   -1203417    +767378
      WHEN 1672 => Ti := "000100111001011100111100110101100010110111101100"; --   +1283900   -2740756
      WHEN 1673 => Ti := "111011010101011111110010000111111110101011011000"; --   -1222670   +2091736
      WHEN 1674 => Ti := "000110000010100000100100000101110001100111010110"; --   +1583140   +1513942
      WHEN 1675 => Ti := "001011101010001111011110111100101110001101100101"; --   +3056606    -859291
      WHEN 1676 => Ti := "110011101010000011010011000011111111110000010010"; --   -3235629   +1047570
      WHEN 1677 => Ti := "110110000011111101110011111111110111011110110000"; --   -2605197     -34896
      WHEN 1678 => Ti := "000000101111011000001100111011010100010011011101"; --    +194060   -1227555
      WHEN 1679 => Ti := "111111110101000100101010001000010100110001111010"; --     -44758   +2182266
      WHEN 1680 => Ti := "000100001111101001100000110111011101010101001101"; --   +1112672   -2239155
      WHEN 1681 => Ti := "110100000000000110101000111100011110110011111000"; --   -3145304    -922376
      WHEN 1682 => Ti := "110100100101101101010000110110001111111011001001"; --   -2991280   -2556215
      WHEN 1683 => Ti := "000001001101001000010111000010111011111111111001"; --    +315927    +770041
      WHEN 1684 => Ti := "000111001101001010100111110111110010001110111011"; --   +1888935   -2153541
      WHEN 1685 => Ti := "110101100000000111001100000000101011000101011100"; --   -2752052    +176476
      WHEN 1686 => Ti := "000100111010011100111101110100011011011010011110"; --   +1287997   -3033442
      WHEN 1687 => Ti := "001001000111110100111011111000101011101111010001"; --   +2391355   -1917999
      WHEN 1688 => Ti := "001010010111101110111111001100101010101101001000"; --   +2718655   +3320648
      WHEN 1689 => Ti := "110101100111001010011100110100010000011010011010"; --   -2723172   -3078502
      WHEN 1690 => Ti := "111000100011111110101111000110110011100100100010"; --   -1949777   +1784098
      WHEN 1691 => Ti := "001010010001010010001010110100101100110000111110"; --   +2692234   -2962370
      WHEN 1692 => Ti := "111111101111100111110101001000001000100001110101"; --     -67083   +2132085
      WHEN 1693 => Ti := "111011011000110011000000111100000111100000100011"; --   -1209152   -1017821
      WHEN 1694 => Ti := "001000110100110001100111000011111010101001110110"; --   +2313319   +1026678
      WHEN 1695 => Ti := "000011100101110010110110111010110101101001101011"; --    +941238   -1353109
      WHEN 1696 => Ti := "000001001101100001111101000001000011101000110010"; --    +317565    +277042
      WHEN 1697 => Ti := "111011001011101111101110111011111001100110110111"; --   -1262610   -1074761
      WHEN 1698 => Ti := "000000010011100001101000111101100101110111100000"; --     +79976    -631328
      WHEN 1699 => Ti := "111100110001111101000111110111110001001000100001"; --    -843961   -2158047
      WHEN 1700 => Ti := "111101110101010111000111110111001111111110101110"; --    -567865   -2293842
      WHEN 1701 => Ti := "000111111101100100011111110100100001001101101101"; --   +2087199   -3009683
      WHEN 1702 => Ti := "110110101001010100011011111001110110100010111001"; --   -2452197   -1611591
      WHEN 1703 => Ti := "000101111111010110111101110100010001010100000000"; --   +1570237   -3074816
      WHEN 1704 => Ti := "000011111100111111110010000111100100010100110100"; --   +1036274   +1983796
      WHEN 1705 => Ti := "000111110010000100011011001100010000011001110010"; --   +2040091   +3212914
      WHEN 1706 => Ti := "110101110100000100000111001000100111000101001101"; --   -2670329   +2257229
      WHEN 1707 => Ti := "000111100001010001001000001011101111111100110010"; --   +1971272   +3079986
      WHEN 1708 => Ti := "110100111000100110111101111100110011010000110011"; --   -2913859    -838605
      WHEN 1709 => Ti := "000101000111010000001110110011101001100011110010"; --   +1340430   -3237646
      WHEN 1710 => Ti := "001001000000010001101011000010111101110011000110"; --   +2360427    +777414
      WHEN 1711 => Ti := "111011000111111001010011001100010100001001110011"; --   -1278381   +3228275
      WHEN 1712 => Ti := "001000101000010100101111001010001100000010100110"; --   +2262319   +2670758
      WHEN 1713 => Ti := "000011010100101100010110110100000001000000101110"; --    +871190   -3141586
      WHEN 1714 => Ti := "000001111100000010001111110100000111000011111101"; --    +508047   -3116803
      WHEN 1715 => Ti := "110101010011111010010100110011101100100011110011"; --   -2802028   -3225357
      WHEN 1716 => Ti := "000111111101011010111001111100010011001010001110"; --   +2086585    -970098
      WHEN 1717 => Ti := "001001100101011110101101110100010101000000110101"; --   +2512813   -3059659
      WHEN 1718 => Ti := "110100100100010000011100111000101000010010011100"; --   -2997220   -1932132
      WHEN 1719 => Ti := "111110101001010100001110111100001001010110111101"; --    -355058   -1010243
      WHEN 1720 => Ti := "001001101110100101001010111001111101000010111100"; --   +2550090   -1584964
      WHEN 1721 => Ti := "111101110001100000101100110100100001110100000111"; --    -583636   -3007225
      WHEN 1722 => Ti := "000010110001011111010110111010100110000110011000"; --    +726998   -1416808
      WHEN 1723 => Ti := "001001110101110001111111000110000111111010101011"; --   +2579583   +1605291
      WHEN 1724 => Ti := "000000001010011110011000001000010011101110101101"; --     +42904   +2177965
      WHEN 1725 => Ti := "000010100100011000111000111111001110010100111010"; --    +673336    -203462
      WHEN 1726 => Ti := "111000000011111011010110111101101011000001001000"; --   -2081066    -610232
      WHEN 1727 => Ti := "000110101010010100000000111000011001110010010111"; --   +1746176   -1991529
      WHEN 1728 => Ti := "111100100101000011011100000101010110110111001100"; --    -896804   +1404364
      WHEN 1729 => Ti := "001011111100111001001100111000001011111011111000"; --   +3133004   -2048264
      WHEN 1730 => Ti := "000010000100011000101100111011001101101101000000"; --    +542252   -1254592
      WHEN 1731 => Ti := "111000000001110100111100111100111110110100000100"; --   -2089668    -791292
      WHEN 1732 => Ti := "110110010000100111011110111111001111010100111011"; --   -2553378    -199365
      WHEN 1733 => Ti := "110110111001110111101110111010110110110000000101"; --   -2384402   -1348603
      WHEN 1734 => Ti := "000101110110111101010011000001100100010101110001"; --   +1535827    +410993
      WHEN 1735 => Ti := "110011101110000011010101000001001010100101101000"; --   -3219243    +305512
      WHEN 1736 => Ti := "111010111110001111101001000001111011101111100001"; --   -1317911    +506849
      WHEN 1737 => Ti := "001010101110001000101110111100000010001101010100"; --   +2810414   -1039532
      WHEN 1738 => Ti := "111000011010111011011111111100111101111101101011"; --   -1986849    -794773
      WHEN 1739 => Ti := "001011101010011001000101111000111000010010100010"; --   +3057221   -1866590
      WHEN 1740 => Ti := "111100010000100110100001110100111101001101110111"; --    -980575   -2894985
      WHEN 1741 => Ti := "111101011111000110111111111011100101111101001010"; --    -659009   -1155254
      WHEN 1742 => Ti := "000111001011100001000000110110110101111000001011"; --   +1882176   -2400757
      WHEN 1743 => Ti := "000111001110110111011011111110110000111110010110"; --   +1895899    -323690
      WHEN 1744 => Ti := "000110010110000000101100001001000100101011110010"; --   +1663020   +2378482
      WHEN 1745 => Ti := "111011110011000011001001111001010111011100010100"; --   -1101623   -1738988
      WHEN 1746 => Ti := "110110111000001110000111111110101101010100101110"; --   -2391161    -338642
      WHEN 1747 => Ti := "000110001010100011110100000100010001101101001100"; --   +1616116   +1121100
      WHEN 1748 => Ti := "111010001110001000111101000010110001101100101000"; --   -1514947    +727848
      WHEN 1749 => Ti := "000000011101000001101011111010000011100110001011"; --    +118891   -1558133
      WHEN 1750 => Ti := "000101101100101101001111001001011110010010010101"; --   +1493839   +2483349
      WHEN 1751 => Ti := "110011011100100000000001111000001011101111000101"; --   -3291135   -2049083
      WHEN 1752 => Ti := "111110001011000111001111111011001101100000001101"; --    -478769   -1255411
      WHEN 1753 => Ti := "111100001001101100111000000010100001110110001000"; --   -1008840    +662920
      WHEN 1754 => Ti := "000011101111011001010100111010010101010110010010"; --    +980564   -1485422
      WHEN 1755 => Ti := "111011011010101100100111111101000100110111010100"; --   -1201369    -766508
      WHEN 1756 => Ti := "001011000011101000110110111101110110111010110011"; --   +2898486    -561485
      WHEN 1757 => Ti := "000000011001011011010000001001100000111111001001"; --    +104144   +2494409
      WHEN 1758 => Ti := "001000010101101011000010001000011110111011100100"; --   +2185922   +2223844
      WHEN 1759 => Ti := "000101000100011101000000111100101001111010010110"; --   +1328960    -876906
      WHEN 1760 => Ti := "111100110011010000010101000011000010100011001000"; --    -838635    +796872
      WHEN 1761 => Ti := "000111001100101010100111111001010011111111100000"; --   +1886887   -1753120
      WHEN 1762 => Ti := "110111010110011011000101000001100110010010100101"; --   -2267451    +418981
      WHEN 1763 => Ti := "111011010110010010111111111110001111001110001001"; --   -1219393    -461943
      WHEN 1764 => Ti := "001100100001011111110011111010011010101001100001"; --   +3282931   -1463711
      WHEN 1765 => Ti := "001010110000101111001001110100101011111010100100"; --   +2821065   -2965852
      WHEN 1766 => Ti := "001001101010111011100010000010101111111111110100"; --   +2535138    +720884
      WHEN 1767 => Ti := "000000000011011110010101110011101010000110111111"; --     +14229   -3235393
      WHEN 1768 => Ti := "000001000000101000010010111111000110000001101010"; --    +264722    -237462
      WHEN 1769 => Ti := "000110110011010000110111111000100100001100000001"; --   +1782839   -1948927
      WHEN 1770 => Ti := "001100000111001001010000110100011111111010100000"; --   +3174992   -3015008
      WHEN 1771 => Ti := "001000010101101011000010111100100100010011111011"; --   +2185922    -899845
      WHEN 1772 => Ti := "111100000010000000000010000010000111011001001011"; --   -1040382    +554571
      WHEN 1773 => Ti := "111101000010000110110100110100001001001010010111"; --    -777804   -3108201
      WHEN 1774 => Ti := "000111111010110001010001111101011001100001000010"; --   +2075729    -681918
      WHEN 1775 => Ti := "111100011001110110100101000110100001110111101000"; --    -942683   +1711592
      WHEN 1776 => Ti := "111110000010001101100101000100111101110000101001"; --    -515227   +1301545
      WHEN 1777 => Ti := "111100111000001101001010001010100101010101111101"; --    -818358   +2774397
      WHEN 1778 => Ti := "001000000100001110001000000100011111011010000100"; --   +2114440   +1177220
      WHEN 1779 => Ti := "110100000000110000001111111101000111110111010101"; --   -3142641    -754219
      WHEN 1780 => Ti := "000110101001010000110011111101101010101010101110"; --   +1741875    -611666
      WHEN 1781 => Ti := "111011001010000110000111111110010011100001010111"; --   -1269369    -444329
      WHEN 1782 => Ti := "111011010110101001011000110111000000010101000010"; --   -1217960   -2357950
      WHEN 1783 => Ti := "110110001011000111011100001010000011000010100011"; --   -2575908   +2633891
      WHEN 1784 => Ti := "000101001010011001110110111110000101101010111001"; --   +1353334    -501063
      WHEN 1785 => Ti := "111001110010111111001101111001000110101100001110"; --   -1626163   -1807602
      WHEN 1786 => Ti := "000000000111010001100011000100011110001010000100"; --     +29795   +1172100
      WHEN 1787 => Ti := "001000110110101011001110111110110011110111111101"; --   +2321102    -311811
      WHEN 1788 => Ti := "111111011110000100100001000100110101100000100110"; --    -138975   +1267750
      WHEN 1789 => Ti := "111111100001100111110000111101110101101010110011"; --    -124432    -566605
      WHEN 1790 => Ti := "111111111001101011000101000100011001011101001111"; --     -25915   +1152847
      WHEN 1791 => Ti := "110111000100010001011000000001101001001100001101"; --   -2341800    +430861
      WHEN 1792 => Ti := "001000111011010100110110110111110000001110111010"; --   +2340150   -2161734
      WHEN 1793 => Ti := "111001001011000101010111000011101110101100111111"; --   -1789609    +977727
      WHEN 1794 => Ti := "000001100110100101010100000101100101110111010010"; --    +420180   +1465810
      WHEN 1795 => Ti := "000000100101101011010101111101100101100100010011"; --    +154325    -632557
      WHEN 1796 => Ti := "001001010001001110100101111011001110111001110100"; --   +2429861   -1249676
      WHEN 1797 => Ti := "000100100100111100110101001000000100001110100111"; --   +1199925   +2114471
      WHEN 1798 => Ti := "111110101110110100010000000111000011000111110101"; --    -332528   +1847797
      WHEN 1799 => Ti := "110011001111001100101111001001000000001011110000"; --   -3345617   +2360048
      WHEN 1800 => Ti := "000110101101100111001110001100101100111001111100"; --   +1759694   +3329660
      WHEN 1801 => Ti := "001011011110011001000000111100101100110011111110"; --   +3008064    -865026
      WHEN 1802 => Ti := "001000101110110100110010110100000011010111001000"; --   +2288946   -3131960
      WHEN 1803 => Ti := "111010100110001001000110110101101010001110001000"; --   -1416634   -2710648
      WHEN 1804 => Ti := "110011001111111100110000111001111011000110001000"; --   -3342544   -1592952
      WHEN 1805 => Ti := "111011001101000010111011111001110000001111101010"; --   -1257285   -1637398
      WHEN 1806 => Ti := "001011000100011111010000111101000101010111010100"; --   +2901968    -764460
      WHEN 1807 => Ti := "001100011111011111110010001010011101001001000110"; --   +3274738   +2740806
      WHEN 1808 => Ti := "111101001001111101010000000001111010100010101101"; --    -745648    +501933
      WHEN 1809 => Ti := "111111100111010001011000111111010011111110100011"; --    -101288    -180317
      WHEN 1810 => Ti := "110110111100011010111100000000101101010010010000"; --   -2373956    +185488
      WHEN 1811 => Ti := "001011111010000101111110000000010010011011101100"; --   +3121534     +75500
      WHEN 1812 => Ti := "111100010001101001101111000101110100100111010111"; --    -976273   +1526231
      WHEN 1813 => Ti := "110100010110010000010111111010010100110011000101"; --   -3054569   -1487675
      WHEN 1814 => Ti := "001011110010010010101110000100011110110110110111"; --   +3089582   +1174967
      WHEN 1815 => Ti := "001000101011011110010111110101011000011010110101"; --   +2275223   -2783563
      WHEN 1816 => Ti := "111100001001000000000101111101000010010000111001"; --   -1011707    -777159
      WHEN 1817 => Ti := "001100100011111100100111001100101101011101001001"; --   +3292967   +3331913
      WHEN 1818 => Ti := "001001010110000001110100001010101001111100011000"; --   +2449524   +2793240
      WHEN 1819 => Ti := "000010011001011100000000001010001011010010100110"; --    +628480   +2667686
      WHEN 1820 => Ti := "111100011101001001110011111001010010011001000110"; --    -929165   -1759674
      WHEN 1821 => Ti := "111101110011010011111010111111000011000001101001"; --    -576262    -249751
      WHEN 1822 => Ti := "111110100110100100001101110111110111011000100011"; --    -366323   -2132445
      WHEN 1823 => Ti := "111011010011100010111110110100100111100000111100"; --   -1230658   -2983876
      WHEN 1824 => Ti := "000001100110101011101101000111100011010100110100"; --    +420589   +1979700
      WHEN 1825 => Ti := "111010111011011111101000110101011111000100011110"; --   -1329176   -2756322
      WHEN 1826 => Ti := "000010010001011111001010001000110110001000100000"; --    +595914   +2318880
      WHEN 1827 => Ti := "110100110011000011101110001001111000011000111001"; --   -2936594   +2590265
      WHEN 1828 => Ti := "110101001001011101011101000111010101101011001000"; --   -2844835   +1923784
      WHEN 1829 => Ti := "111111000000010001001010000001011100001100001000"; --    -261046    +377608
      WHEN 1830 => Ti := "001000000110000100100010001011010100000110001110"; --   +2122018   +2965902
      WHEN 1831 => Ti := "001000101110011110011000001011001111101100100110"; --   +2287512   +2947878
      WHEN 1832 => Ti := "001001100001111110101011111000011001100101100011"; --   +2498475   -1992349
      WHEN 1833 => Ti := "000001110010011110111110110110011111001000000010"; --    +468926   -2493950
      WHEN 1834 => Ti := "000110001000100000100111110011101011011101011001"; --   +1607719   -3229863
      WHEN 1835 => Ti := "000101111000110110111010000011000000101001100001"; --   +1543610    +789089
      WHEN 1836 => Ti := "000111010111100001000100001011101000100110010110"; --   +1931332   +3049878
      WHEN 1837 => Ti := "111100001111111001101110000010011110010010111010"; --    -983442    +648378
      WHEN 1838 => Ti := "000011101011101100011111000010101111111100100111"; --    +965407    +720679
      WHEN 1839 => Ti := "110110001001000100001111111110001100010001010101"; --   -2584305    -474027
      WHEN 1840 => Ti := "000100010110101100101111110111001010111011100000"; --   +1141551   -2314528
      WHEN 1841 => Ti := "001001110110101011100110001000110011101110111001"; --   +2583270   +2309049
      WHEN 1842 => Ti := "111000001010101110100110111011011010010000010010"; --   -2053210   -1203182
      WHEN 1843 => Ti := "110100011111101010000001001001011010111111000111"; --   -3016063   +2469831
      WHEN 1844 => Ti := "000011110001001100100001110100000101100111001001"; --    +987937   -3122743
      WHEN 1845 => Ti := "110011011110010110011100110100001010100011111110"; --   -3283556   -3102466
      WHEN 1846 => Ti := "111010000010100101101100000001111100101100010100"; --   -1562260    +510740
      WHEN 1847 => Ti := "000110011010010000101101001010101001001111100101"; --   +1680429   +2790373
      WHEN 1848 => Ti := "000000100011111011010100111111010011010100111100"; --    +147156    -182980
      WHEN 1849 => Ti := "001010010010101000100100111110100101110100101011"; --   +2697764    -369365
      WHEN 1850 => Ti := "001010011110101111000010001011010101100110001111"; --   +2747330   +2972047
      WHEN 1851 => Ti := "111000010011001000001111110111100111101011101010"; --   -2018801   -2196758
      WHEN 1852 => Ti := "111010101010011100010101110111010001000001111011"; --   -1399019   -2289541
      WHEN 1853 => Ti := "000101111000001010000111001001100101101111001011"; --   +1540743   +2513867
      WHEN 1854 => Ti := "111101111001000000101111110110001000110100101101"; --    -552913   -2585299
      WHEN 1855 => Ti := "001010000010001000011110000010110101001001011100"; --   +2630174    +741980
      WHEN 1856 => Ti := "000111011111001010101101111100111000010111001111"; --   +1962669    -817713
      WHEN 1857 => Ti := "111111000111011010110011000110001110111010101110"; --    -231757   +1633966
      WHEN 1858 => Ti := "000001001101100101001010000000001101011000011110"; --    +317770     +54814
      WHEN 1859 => Ti := "000101000001111001110011001011100100010011000111"; --   +1318515   +3032263
      WHEN 1860 => Ti := "111111001101101110000010111101111110110001010000"; --    -205950    -529328
      WHEN 1861 => Ti := "000111111001001110000100000110110111000111110000"; --   +2069380   +1798640
      WHEN 1862 => Ti := "001000110011101011001101111111100110000001110110"; --   +2308813    -106378
      WHEN 1863 => Ti := "001000110000111011001100000100011011111010000011"; --   +2297548   +1162883
      WHEN 1864 => Ti := "111010000111010010100001000011000010111100101110"; --   -1543007    +798510
      WHEN 1865 => Ti := "111001001100100010001011111010011000000110010011"; --   -1783669   -1474157
      WHEN 1866 => Ti := "110101110000111010011111111000001110101011111001"; --   -2683233   -2036999
      WHEN 1867 => Ti := "110100000011111101000011000011011101110000000101"; --   -3129533    +908293
      WHEN 1868 => Ti := "000100001110101100101100001100111001010011100111"; --   +1108780   +3380455
      WHEN 1869 => Ti := "110111100111011011001100110111100011001011101001"; --   -2197812   -2215191
      WHEN 1870 => Ti := "001011001101011100000111110100110101110100001110"; --   +2938631   -2925298
      WHEN 1871 => Ti := "000100110011101100111010111011110010100110110101"; --   +1260346   -1103435
      WHEN 1872 => Ti := "000111011110110111100001000010011000101100011111"; --   +1961441    +625439
      WHEN 1873 => Ti := "111011000011000010110111111110101101111011001000"; --   -1298249    -336184
      WHEN 1874 => Ti := "000000011000101110011101001001011100101111001000"; --    +101277   +2477000
      WHEN 1875 => Ti := "111010110101000101111111000111010111110111111101"; --   -1355393   +1932797
      WHEN 1876 => Ti := "000101110001010000011110111010111010110110100000"; --   +1512478   -1331808
      WHEN 1877 => Ti := "110011001011111111111011111110101011011110010100"; --   -3358725    -346220
      WHEN 1878 => Ti := "111100010111110011010111111111011101001110100110"; --    -951081    -142426
      WHEN 1879 => Ti := "001010110100011000110001110011111000001010010001"; --   +2836017   -3177839
      WHEN 1880 => Ti := "001001011110001110101010111111010101101000001010"; --   +2483114    -173558
      WHEN 1881 => Ti := "001000110101101011001110000011001100110110011001"; --   +2317006    +839065
      WHEN 1882 => Ti := "111011010111110010111111111000001010100101011110"; --   -1213249   -2053794
      WHEN 1883 => Ti := "000111100111000100010111111001001100100010101010"; --   +1995031   -1783638
      WHEN 1884 => Ti := "111111100010110100100011110100011010111010011110"; --    -119517   -3035490
      WHEN 1885 => Ti := "111100000000000000000010110011100000110110111011"; --   -1048574   -3273285
      WHEN 1886 => Ti := "000100000001001001011010000101101010100111010100"; --   +1053274   +1485268
      WHEN 1887 => Ti := "110101000110010000101001111111111011011110110010"; --   -2857943     -18510
      WHEN 1888 => Ti := "111011001110000110001000111011110010101010000010"; --   -1252984   -1103230
      WHEN 1889 => Ti := "000101001011101001110110111010011010110011000111"; --   +1358454   -1463097
      WHEN 1890 => Ti := "111001011110000101011110000110111011110100100101"; --   -1711778   +1817893
      WHEN 1891 => Ti := "000100101110110000000101110111111001001110111110"; --   +1240069   -2124866
      WHEN 1892 => Ti := "111100111010100000010111111110011010010111110100"; --    -808937    -416268
      WHEN 1893 => Ti := "000110101100011010011010111110011000001011000000"; --   +1754778    -425280
      WHEN 1894 => Ti := "001010010100011110111110111010010101111001011111"; --   +2705342   -1483169
      WHEN 1895 => Ti := "111011100110100110010010001011011011011001011110"; --   -1152622   +2995806
      WHEN 1896 => Ti := "001001000111011000001000111010010010001111110111"; --   +2389512   -1498121
      WHEN 1897 => Ti := "110100010110000110110000110110011010101110011010"; --   -3055184   -2511974
      WHEN 1898 => Ti := "001001000101001011010100111001110000000110000100"; --   +2380500   -1638012
      WHEN 1899 => Ti := "000010001010111011111011111100010001100000100111"; --    +569083    -976857
      WHEN 1900 => Ti := "110101101100000100000100111001110000010110000100"; --   -2703100   -1636988
      WHEN 1901 => Ti := "001011001010001100000101000010001111001100011011"; --   +2925317    +586523
      WHEN 1902 => Ti := "111011000110010010111001111001110100000110000101"; --   -1284935   -1621627
      WHEN 1903 => Ti := "110111001000101110001101110110111001101011011001"; --   -2323571   -2385191
      WHEN 1904 => Ti := "000111001011111101110011000001001101001111001111"; --   +1884019    +316367
      WHEN 1905 => Ti := "001100001111111100100000111000101100010101101010"; --   +3211040   -1915542
      WHEN 1906 => Ti := "110111011100100100101110111111101011000001111000"; --   -2242258     -85896
      WHEN 1907 => Ti := "111000110000101000011010110101110010100100100101"; --   -1897958   -2676443
      WHEN 1908 => Ti := "110111101110101011001110001100110001000000010111"; --   -2168114   +3346455
      WHEN 1909 => Ti := "111010111011111111101000000110010100000100010110"; --   -1327128   +1655062
      WHEN 1910 => Ti := "001001000001111000000110000000010000011110111000"; --   +2366982     +67512
      WHEN 1911 => Ti := "001010111101000010011010000001100010011100001010"; --   +2871450    +403210
      WHEN 1912 => Ti := "000001000111111000010101000100011001010000011100"; --    +294421   +1152028
      WHEN 1913 => Ti := "110111101001101110011001110101011000101110000010"; --   -2188391   -2782334
      WHEN 1914 => Ti := "111010010001010010100101000010110010110110001111"; --   -1502043    +732559
      WHEN 1915 => Ti := "110011110001101100111100000000111101000010010110"; --   -3204292    +250006
      WHEN 1916 => Ti := "000011101111110010111010001100110011011001111111"; --    +982202   +3356287
      WHEN 1917 => Ti := "000100011011000011001010000110000100110100010001"; --   +1159370   +1592593
      WHEN 1918 => Ti := "001010011011101111000001000110011111110100011011"; --   +2735041   +1703195
      WHEN 1919 => Ti := "000001100011011110111001111111100100001011011100"; --    +407481    -113956
      WHEN 1920 => Ti := "111101011101010110111110000001111011111001000111"; --    -666178    +507463
      WHEN 1921 => Ti := "111111110001110001011100001001101100100101100111"; --     -58276   +2541927
      WHEN 1922 => Ti := "001100011111111100100110111000010001001011111010"; --   +3276582   -2026758
      WHEN 1923 => Ti := "000111010110100100010001000100000111100000010101"; --   +1927441   +1079317
      WHEN 1924 => Ti := "000011101100101111101100000001011110111000111100"; --    +969708    +388668
      WHEN 1925 => Ti := "001001010000010100111110110100011100001010011110"; --   +2426174   -3030370
      WHEN 1926 => Ti := "001001010010000100111111000101001101010011111100"; --   +2433343   +1365244
      WHEN 1927 => Ti := "110110010010110111011111110111000100010001110111"; --   -2544161   -2341769
      WHEN 1928 => Ti := "110011111110101001110100000101010111101101100110"; --   -3151244   +1407846
      WHEN 1929 => Ti := "000010101100000101101110111111000100000001101010"; --    +704878    -245654
      WHEN 1930 => Ti := "111110010100110111010011111101000110001101101110"; --    -438829    -760978
      WHEN 1931 => Ti := "111010000011111100000110111111011111011000001101"; --   -1556730    -133619
      WHEN 1932 => Ti := "110100011001010011100101110100101010101101110000"; --   -3042075   -2970768
      WHEN 1933 => Ti := "111011000111111001010011001011110010001001100110"; --   -1278381   +3088998
      WHEN 1934 => Ti := "000110011001101010010011111000000111011000101001"; --   +1677971   -2066903
      WHEN 1935 => Ti := "111110111110110001001001001001100100111000110001"; --    -267191   +2510385
      WHEN 1936 => Ti := "110111010100011011000101110111101011110101010010"; --   -2275643   -2179758
      WHEN 1937 => Ti := "000011010011011001001001000001100101011000111111"; --    +865865    +415295
      WHEN 1938 => Ti := "000101001101000000010000001100100010000011011111"; --   +1363984   +3285215
      WHEN 1939 => Ti := "001000001000110001010111110110101110100100111011"; --   +2133079   -2430661
      WHEN 1940 => Ti := "110101011111111101100110110101101010111110001000"; --   -2752666   -2707576
      WHEN 1941 => Ti := "000101010111111001111011000100010100011010000000"; --   +1408635   +1132160
      WHEN 1942 => Ti := "001001011101100001110110111010110011000110011101"; --   +2480246   -1363555
      WHEN 1943 => Ti := "001000101010100100110000110111010001010101001000"; --   +2271536   -2288312
      WHEN 1944 => Ti := "111000001010100001110010001000111010111011101110"; --   -2054030   +2338542
      WHEN 1945 => Ti := "000110001011111010001110001001100110100101100101"; --   +1621646   +2517349
      WHEN 1946 => Ti := "111111000001101010110000000011010001010000000001"; --    -255312    +857089
      WHEN 1947 => Ti := "110011011101000000000001110100001000111101100100"; --   -3289087   -3109020
      WHEN 1948 => Ti := "110011000111101001100000000010110110111111110111"; --   -3376544    +749559
      WHEN 1949 => Ti := "000011011001001100011000111101101101111010110000"; --    +889624    -598352
      WHEN 1950 => Ti := "111101110010001010010011111111000101001011010000"; --    -580973    -240944
      WHEN 1951 => Ti := "000001001111111011100101001000100101101011100110"; --    +327397   +2251494
      WHEN 1952 => Ti := "001000011100111011000101000000001010011000011100"; --   +2215621     +42524
      WHEN 1953 => Ti := "000111111101000100011111111000100000110010011001"; --   +2085151   -1962855
      WHEN 1954 => Ti := "000010001001001111000111001001000100001011110010"; --    +562119   +2376434
      WHEN 1955 => Ti := "111001111100011000110111001011111000100011001111"; --   -1587657   +3115215
      WHEN 1956 => Ti := "000010100111100010011111001100110101111010000000"; --    +686239   +3366528
      WHEN 1957 => Ti := "110111000001100111110001000010010011001111101001"; --   -2352655    +603113
      WHEN 1958 => Ti := "110101100010110100000000000011011100000110011110"; --   -2740992    +901534
      WHEN 1959 => Ti := "000001000101101110101110110111110011101000100010"; --    +285614   -2147806
      WHEN 1960 => Ti := "000100111101100011010111001011100011001111111010"; --   +1300695   +3027962
      WHEN 1961 => Ti := "110011101011000011010100000010010111000010111000"; --   -3231532    +618680
      WHEN 1962 => Ti := "000110111101000100000111111010010100001100101011"; --   +1822983   -1490133
      WHEN 1963 => Ti := "111111001011110111100111111000110000101100000110"; --    -213529   -1897722
      WHEN 1964 => Ti := "001100001100111001010010111001101011100110000010"; --   +3198546   -1656446
      WHEN 1965 => Ti := "111110111101100111100010001010001111001100001110"; --    -271902   +2683662
      WHEN 1966 => Ti := "000110100100001101100100111100100110001101100010"; --   +1721188    -892062
      WHEN 1967 => Ti := "110100100101101010000011110100010000100111001101"; --   -2991485   -3077683
      WHEN 1968 => Ti := "001011101110111100010011110110101010111011010100"; --   +3075859   -2445612
      WHEN 1969 => Ti := "111111101010010111110011111101110101101010110011"; --     -88589    -566605
      WHEN 1970 => Ti := "110111111001101110011111000100111000000000100111"; --   -2122849   +1277991
      WHEN 1971 => Ti := "000010110011101100001010000101110101011101110001"; --    +736010   +1529713
      WHEN 1972 => Ti := "110100100001111010000010110100111001001010101001"; --   -3006846   -2911575
      WHEN 1973 => Ti := "000000010110000001101001111110101111100111111011"; --     +90217    -329221
      WHEN 1974 => Ti := "110011111010100110100110001011111011110000000011"; --   -3167834   +3128323
      WHEN 1975 => Ti := "111001000000000101010011001011111011100110011101"; --   -1834669   +3127709
      WHEN 1976 => Ti := "001100000011001100011011111010100100001001100100"; --   +3158811   -1424796
      WHEN 1977 => Ti := "001010010010010101010111000001000110000010011001"; --   +2696535    +286873
      WHEN 1978 => Ti := "110100101100000000011111111000000010101011110100"; --   -2965473   -2086156
      WHEN 1979 => Ti := "111101010010011010000111111000000000100010001101"; --    -711033   -2094963
      WHEN 1980 => Ti := "111001100001000101100000001100001111100011011000"; --   -1699488   +3209432
      WHEN 1981 => Ti := "000011100100000010110110001010000110001000111110"; --    +934070   +2646590
      WHEN 1982 => Ti := "001010101110011000101110000010101010111001011001"; --   +2811438    +699993
      WHEN 1983 => Ti := "000110000010001010001011111011011100101001111001"; --   +1581707   -1193351
      WHEN 1984 => Ti := "001001101001011000010100110100000111100111001010"; --   +2528788   -3114550
      WHEN 1985 => Ti := "110110110000100001010001111110100001001110010000"; --   -2422703    -388208
      WHEN 1986 => Ti := "111011110110111100110001111010111110000011010100"; --   -1085647   -1318700
      WHEN 1987 => Ti := "001001100011101011011111110111101000111110111000"; --   +2505439   -2191432
      WHEN 1988 => Ti := "110101100001010000110011111111101111001110101101"; --   -2747341     -68691
      WHEN 1989 => Ti := "110111011101010111111011000001001101001111001111"; --   -2238981    +316367
      WHEN 1990 => Ti := "111110111101010100010101111110101011111011000111"; --    -273131    -344377
      WHEN 1991 => Ti := "111101110101011010010100111110000110001010111001"; --    -567660    -499015
      WHEN 1992 => Ti := "111001100000100010010011000000110111111011111010"; --   -1701741    +229114
      WHEN 1993 => Ti := "001001111100111011101001111011001010001100111111"; --   +2608873   -1268929
      WHEN 1994 => Ti := "111010110011111111100101110110010000010111111101"; --   -1359899   -2554371
      WHEN 1995 => Ti := "110100111111011101011010111010001000110110001101"; --   -2885798   -1536627
      WHEN 1996 => Ti := "001000111100111110011101111000000010111000101000"; --   +2346909   -2085336
      WHEN 1997 => Ti := "110100100001100011101000000000011100101110111101"; --   -3008280    +117693
      WHEN 1998 => Ti := "111011011100010011000001000111010011101011001000"; --   -1194815   +1915592
      WHEN 1999 => Ti := "001001110011111110110010000100001101010011100100"; --   +2572210   +1103076
      WHEN 2000 => Ti := "000101000100101001110100000010001101101111100111"; --   +1329780    +580583
      WHEN 2001 => Ti := "111010011000000010100111111000010011110010010100"; --   -1474393   -2016108
      WHEN 2002 => Ti := "110111011001010001100000111101100011011101111001"; --   -2255776    -641159
      WHEN 2003 => Ti := "000010100111111100000110111000010110111000101111"; --    +687878   -2003409
      WHEN 2004 => Ti := "110111000100011010111111001001101011100010011010"; --   -2341185   +2537626
      WHEN 2005 => Ti := "000000000110100001100011001000011100011000010110"; --     +26723   +2213398
      WHEN 2006 => Ti := "111110101001100100001110110110111010000001110011"; --    -354034   -2383757
      WHEN 2007 => Ti := "110111011010101011000111000011001010011100110001"; --   -2250041    +829233
      WHEN 2008 => Ti := "000000100111110100111100000110111110110100100110"; --    +163132   +1830182
      WHEN 2009 => Ti := "000000001100111110011000110110101101101000001000"; --     +53144   -2434552
      WHEN 2010 => Ti := "000110010011101010010001000101111101101101110100"; --   +1653393   +1563508
      WHEN 2011 => Ti := "111011001000010010111001001011011010001001011101"; --   -1276743   +2990685
      WHEN 2012 => Ti := "000010110010010010100011000101000000000011110111"; --    +730275   +1310967
      WHEN 2013 => Ti := "000010110001111111010110000001010000011000110111"; --    +729046    +329271
      WHEN 2014 => Ti := "000100010011010011001000111110000111010001010011"; --   +1127624    -494509
      WHEN 2015 => Ti := "111011010110101111110010111000100110000010011011"; --   -1217550   -1941349
      WHEN 2016 => Ti := "111011010010110010111101000001110111000101111000"; --   -1233731    +487800
      WHEN 2017 => Ti := "111110110110000100010011111001110000111111101011"; --    -302829   -1634325
      WHEN 2018 => Ti := "110100101100010011101100000010110101011111110110"; --   -2964244    +743414
      WHEN 2019 => Ti := "001001101001000001111011001001011100011000101110"; --   +2527355   +2475566
      WHEN 2020 => Ti := "111110101010001010101000111001011011000010101111"; --    -351576   -1724241
      WHEN 2021 => Ti := "001011100110101100010000001010011010001100010010"; --   +3042064   +2728722
      WHEN 2022 => Ti := "111011110001010110010110110011110011001101011100"; --   -1108586   -3198116
      WHEN 2023 => Ti := "110100110001111101010100000111001011111011000101"; --   -2941100   +1883845
      WHEN 2024 => Ti := "000010010001011000110000111111110010101110101110"; --    +595504     -54354
      WHEN 2025 => Ti := "111011010111101100100110001010101101100110000000"; --   -1213658   +2808192
      WHEN 2026 => Ti := "001011010110101000111101000010100100100010111101"; --   +2976317    +673981
      WHEN 2027 => Ti := "111110111011101010101110001000110111110101010100"; --    -279890   +2325844
      WHEN 2028 => Ti := "110110011111111101111110000101011010010111001110"; --   -2490498   +1418702
      WHEN 2029 => Ti := "111001101010010010010110111110000100100001010010"; --   -1661802    -505774
      WHEN 2030 => Ti := "001011010010001000111100001011011111110011000110"; --   +2957884   +3013830
      WHEN 2031 => Ti := "111101010011000011101101111001110111011001010011"; --    -708371   -1608109
      WHEN 2032 => Ti := "111101100101110011110100110111111101101011110011"; --    -631564   -2106637
      WHEN 2033 => Ti := "111001010010111000100111001000101001010101001110"; --   -1757657   +2266446
      WHEN 2034 => Ti := "000101001000100011011011111110100111100111111001"; --   +1345755    -361991
      WHEN 2035 => Ti := "111011000010010010110111111101001001100111010101"; --   -1301321    -747051
      WHEN 2036 => Ti := "001100001010111001010001001100111000010000011010"; --   +3190353   +3376154
      WHEN 2037 => Ti := "001100000110001100011100110100010000101010011010"; --   +3171100   -3077478
      WHEN 2038 => Ti := "000110010011101010010001001011110001100110011001"; --   +1653393   +3086745
      WHEN 2039 => Ti := "111000111101010101010010111010001110000011000010"; --   -1845934   -1515326
      WHEN 2040 => Ti := "110011010101011111111111000010001101110010110100"; --   -3319809    +580788
      WHEN 2041 => Ti := "001010100101101000101011111000100000101000110011"; --   +2775595   -1963469
      WHEN 2042 => Ti := "000101010101010000010011111000010010000101100001"; --   +1397779   -2023071
      WHEN 2043 => Ti := "111101001110110000011111000110110010011010111011"; --    -725985   +1779387
      WHEN 2044 => Ti := "000111100100111010110000001001001011111000101000"; --   +1986224   +2407976
      WHEN 2045 => Ti := "001011101100101111011111111001001111111111011110"; --   +3066847   -1769506
      WHEN 2046 => Ti := "111101100100010000100111000100101010010011101111"; --    -637913   +1221871
      WHEN 2047 => Ti := "110011000100010011000101111010000100111111110010"; --   -3390267   -1552398
      WHEN OTHERS => NULL;
    END CASE; 
    T <= Ti; 
  END PROCESS; 
END ARCHITECTURE arch_rom; 



-----------------------------------------------------------
LIBRARY IEEE; 
  USE IEEE.std_logic_1164.all; 

ENTITY goldvect2 IS 
  PORT ( 
    A : IN integer; 
    T : OUT std_logic_vector(47 DOWNTO 0));
END ENTITY goldvect2; 

ARCHITECTURE arch_rom OF goldvect2 IS 
BEGIN 
  PROCESS (A) 
    VARIABLE Ti  : std_logic_vector(47 DOWNTO 0); 
  BEGIN 
    CASE A IS  
      WHEN    0 => Ti := "111111111111111111110110111111111111111111110011"; --        -10        -13
      WHEN    1 => Ti := "000000100101010100110101111011001001001001101001"; --    +152885   -1273239
      WHEN    2 => Ti := "000000000011001101101110000010100101111001001111"; --     +13166    +679503
      WHEN    3 => Ti := "111110100000101001111111111101110011010111111010"; --    -390529    -576006
      WHEN    4 => Ti := "111101110110100110010111000111010011000101101110"; --    -562793   +1913198
      WHEN    5 => Ti := "111100111110101001101010111111001101011010011001"; --    -791958    -207207
      WHEN    6 => Ti := "111111110110110011010000000001101111100101100011"; --     -37680    +457059
      WHEN    7 => Ti := "111111001100101010010011111100100111000011101110"; --    -210285    -888594
      WHEN    8 => Ti := "111110101000100110111110000000001100100110000011"; --    -357954     +51587
      WHEN    9 => Ti := "111110001111001010010000000011000100100101010111"; --    -462192    +805207
      WHEN   10 => Ti := "000001010010100010111111000000110010010001100010"; --    +338111    +205922
      WHEN   11 => Ti := "000010111110010100001111111101100001100010010111"; --    +779535    -649065
      WHEN   12 => Ti := "000011101010000110011001111111110000011001110100"; --    +958873     -63884
      WHEN   13 => Ti := "111110000011011001100101111111000101110110010011"; --    -510363    -238189
      WHEN   14 => Ti := "111110100000010101011010111101001000001011011110"; --    -391846    -752930
      WHEN   15 => Ti := "000000011011001010011100000001001101111101011001"; --    +111260    +319321
      WHEN   16 => Ti := "000000100101100101110011000001100000110110001000"; --    +153971    +396680
      WHEN   17 => Ti := "000011001111011110011101111111010000101111001110"; --    +849821    -193586
      WHEN   18 => Ti := "111100000101010100101111000010100011110000010010"; --   -1026769    +670738
      WHEN   19 => Ti := "000000100111110001011111000001101011101010000110"; --    +162911    +440966
      WHEN   20 => Ti := "000001011110011010011010111110000001000111001111"; --    +386714    -519729
      WHEN   21 => Ti := "111111000001000100000010000010001010100011101001"; --    -257790    +567529
      WHEN   22 => Ti := "000011001111111001111111111100111010110100111010"; --    +851583    -807622
      WHEN   23 => Ti := "000010000000001100010000111110111110101111011001"; --    +525072    -267303
      WHEN   24 => Ti := "000000011000000000000100111101110010000000010111"; --     +98308    -581609
      WHEN   25 => Ti := "111111110010000101001011000001000011000111010011"; --     -57013    +274899
      WHEN   26 => Ti := "000001101011000101101011111100000111001010111111"; --    +438635   -1019201
      WHEN   27 => Ti := "000001101010000100110001111101101110010111001100"; --    +434481    -596532
      WHEN   28 => Ti := "000001111100110010101100111111011000111110110110"; --    +511148    -159818
      WHEN   29 => Ti := "111111101110111001011010000000001110101110000010"; --     -70054     +60290
      WHEN   30 => Ti := "000000111110100000011101000000101011110101101001"; --    +256029    +179561
      WHEN   31 => Ti := "111111010110000110001010111101011111101101110100"; --    -171638    -656524
      WHEN   32 => Ti := "000000010011111000101100000000111000101111001100"; --     +81452    +232396
      WHEN   33 => Ti := "111101111010100001001110111100101111010101101011"; --    -546738    -854677
      WHEN   34 => Ti := "000001100100111110011101111011100010110101010101"; --    +413597   -1168043
      WHEN   35 => Ti := "000010110111100100011000000010000010111010100100"; --    +751896    +536228
      WHEN   36 => Ti := "000100101010000011111001111101010010000010010000"; --   +1220857    -712560
      WHEN   37 => Ti := "000001010111111011001000111111110011010110010010"; --    +360136     -51822
      WHEN   38 => Ti := "111100110100110100101110111101010101111001010001"; --    -832210    -696751
      WHEN   39 => Ti := "111100001101110101001111111100110101110111001100"; --    -991921    -827956
      WHEN   40 => Ti := "000001110100011110011101111111110011010100101101"; --    +477085     -51923
      WHEN   41 => Ti := "111010001111100101101110111110110100100101001100"; --   -1509010    -308916
      WHEN   42 => Ti := "000100010000001001011111111101101011010010001000"; --   +1114719    -609144
      WHEN   43 => Ti := "111110010111010110111001111101111110001110100001"; --    -428615    -531551
      WHEN   44 => Ti := "000001111000000101110101111111110000110000101001"; --    +491893     -62423
      WHEN   45 => Ti := "111111010110110010110101111110111100101111001001"; --    -168779    -275511
      WHEN   46 => Ti := "111110001111111110001000111111000001001010110100"; --    -458872    -257356
      WHEN   47 => Ti := "000100100101010101001000111111010101001010001110"; --   +1201480    -175474
      WHEN   48 => Ti := "111101110001101111011001000010000001110010100101"; --    -582695    +531621
      WHEN   49 => Ti := "000100011001011011111111111111110001011001011011"; --   +1152767     -59813
      WHEN   50 => Ti := "000010100011110000101101000000010000101001001000"; --    +670765     +68168
      WHEN   51 => Ti := "000001001010000111001001111110001010010000010110"; --    +303561    -482282
      WHEN   52 => Ti := "000100111001111000100000111101010101111000110001"; --   +1285664    -696783
      WHEN   53 => Ti := "111010110111000100011000111101000011000010100001"; --   -1347304    -773983
      WHEN   54 => Ti := "000001000110110111101000000010011101011111111111"; --    +290280    +645119
      WHEN   55 => Ti := "000011010100001010001010000010100110011010001100"; --    +869002    +681612
      WHEN   56 => Ti := "111101111111110111111101111111000011001010101111"; --    -524803    -249169
      WHEN   57 => Ti := "111110010110111100010101111111100000101101010001"; --    -430315    -128175
      WHEN   58 => Ti := "000010000010100101010111111101110100111111101111"; --    +534871    -569361
      WHEN   59 => Ti := "000011100101100111010001000000010000100000110001"; --    +940497     +67633
      WHEN   60 => Ti := "000000000110010110010110000100111011010111101100"; --     +26006   +1291756
      WHEN   61 => Ti := "111101001101100111100011000000110001100101101101"; --    -730653    +203117
      WHEN   62 => Ti := "111101110001011010001011000000011110110110100011"; --    -584053    +126371
      WHEN   63 => Ti := "111111111110101011100010000000010011010111001010"; --      -5406     +79306
      WHEN   64 => Ti := "000010001001010100000001111110111010100101110110"; --    +562433    -284298
      WHEN   65 => Ti := "000000101010001000001011000011001111000011110000"; --    +172555    +848112
      WHEN   66 => Ti := "000011110001000001110010111111100110001110110101"; --    +987250    -105547
      WHEN   67 => Ti := "111110110100011001000010111100001010000011111000"; --    -309694   -1007368
      WHEN   68 => Ti := "111111011100010011011110111110100111100111101010"; --    -146210    -362006
      WHEN   69 => Ti := "000001001001010110101011111101010110110111100001"; --    +300459    -692767
      WHEN   70 => Ti := "111110110100101110011111111111000101111000110010"; --    -308321    -238030
      WHEN   71 => Ti := "111101001011111111110001111101011100100000010001"; --    -737295    -669679
      WHEN   72 => Ti := "000011000110100001000011111110111110000000001111"; --    +813123    -270321
      WHEN   73 => Ti := "111111111101000001001010111001010000011011111011"; --     -12214   -1767685
      WHEN   74 => Ti := "000001001011001100100110000010011011001111010000"; --    +308006    +635856
      WHEN   75 => Ti := "111111111001110000110001111110000101001101001000"; --     -25551    -502968
      WHEN   76 => Ti := "000010110000100010011011111101110001001111011010"; --    +723099    -584742
      WHEN   77 => Ti := "111111111000110101111111000001000001000000011010"; --     -29313    +266266
      WHEN   78 => Ti := "111111010000011111001111000100000001011010000000"; --    -194609   +1054336
      WHEN   79 => Ti := "111101111110111011111100111101110011010010000101"; --    -528644    -576379
      WHEN   80 => Ti := "000101110111011111000010111110100011010111001111"; --   +1537986    -379441
      WHEN   81 => Ti := "111101101000100010111001000000110000011100000011"; --    -620359    +198403
      WHEN   82 => Ti := "111100110111000010100100111110111100100010011110"; --    -823132    -276322
      WHEN   83 => Ti := "000100001000111011100000111101111110110011101101"; --   +1085152    -529171
      WHEN   84 => Ti := "111100011101000110001011000001111011100111001010"; --    -929397    +506314
      WHEN   85 => Ti := "000000011100101001100011000100010111101100100100"; --    +117347   +1145636
      WHEN   86 => Ti := "000000001010101001011010000001000111001010110011"; --     +43610    +291507
      WHEN   87 => Ti := "000010011001110001100011111110001001011010000000"; --    +629859    -485760
      WHEN   88 => Ti := "111101010011011110110110111111100110011011110011"; --    -706634    -104717
      WHEN   89 => Ti := "111001011011001001100111000001001010001001100111"; --   -1723801    +303719
      WHEN   90 => Ti := "111110100011011010100110000010100000000110010101"; --    -379226    +655765
      WHEN   91 => Ti := "000010010111100110110011111101110011001111000001"; --    +620979    -576575
      WHEN   92 => Ti := "111110100100001001001110000011011001001101100011"; --    -376242    +889699
      WHEN   93 => Ti := "000001010110101101100000000000100010101111001110"; --    +355168    +142286
      WHEN   94 => Ti := "000001001100000110011111000000001011111011101010"; --    +311711     +48874
      WHEN   95 => Ti := "000110001110110100001001000011001101101101010100"; --   +1633545    +842580
      WHEN   96 => Ti := "000010011001011010100101111101110110010101010100"; --    +628389    -563884
      WHEN   97 => Ti := "000001111101011011110011000000010000001111110110"; --    +513779     +66550
      WHEN   98 => Ti := "000100110101001010111010000001011000000110011010"; --   +1266362    +360858
      WHEN   99 => Ti := "000000100001000101110101111110111110101101110101"; --    +135541    -267403
      WHEN  100 => Ti := "111101111001000100101001111011011000111110101110"; --    -552663   -1208402
      WHEN  101 => Ti := "000000111111010111001110111110000011000001101010"; --    +259534    -511894
      WHEN  102 => Ti := "111101011000010111110000000001000001101100001101"; --    -686608    +269069
      WHEN  103 => Ti := "111111110100110110000001000000001010101100111011"; --     -45695     +43835
      WHEN  104 => Ti := "111011111111110001100010000010111101000101100011"; --   -1049502    +774499
      WHEN  105 => Ti := "111111001001001101011100000000101001000111110011"; --    -224420    +168435
      WHEN  106 => Ti := "111111001001010111100110111111010101111001001111"; --    -223770    -172465
      WHEN  107 => Ti := "000001111011111101000110000010001110001111001110"; --    +507718    +582606
      WHEN  108 => Ti := "111110111101010001110010000010001000000101100100"; --    -273294    +557412
      WHEN  109 => Ti := "111111001110010110001111000000110010011100011001"; --    -203377    +206617
      WHEN  110 => Ti := "000000001010111001111101000010101111110001100111"; --     +44669    +719975
      WHEN  111 => Ti := "111101100011001011100100111100010100001111101110"; --    -642332    -965650
      WHEN  112 => Ti := "111111101000011100001100000001101001101101111111"; --     -96500    +433023
      WHEN  113 => Ti := "111110101001111110011010000010011111100011101100"; --    -352358    +653548
      WHEN  114 => Ti := "000100001011010010011001111111101111110001101011"; --   +1094809     -66453
      WHEN  115 => Ti := "000011101010011000101110000110000001011101111101"; --    +960046   +1578877
      WHEN  116 => Ti := "111111011101100001111000000000101111011111010111"; --    -141192    +194519
      WHEN  117 => Ti := "111110101011111000111111111010100111110011100100"; --    -344513   -1409820
      WHEN  118 => Ti := "000000011101001000011100111110110101000101000000"; --    +119324    -306880
      WHEN  119 => Ti := "111111000111110101101101000000001100010110010101"; --    -230035     +50581
      WHEN  120 => Ti := "111110101101101000101001000011000001110000101111"; --    -337367    +793647
      WHEN  121 => Ti := "000011000110111000111101111101110101100011010100"; --    +814653    -567084
      WHEN  122 => Ti := "000010011010111001000110000001001010010100000110"; --    +634438    +304390
      WHEN  123 => Ti := "000000110010111010001010000000101010110111110010"; --    +208522    +175602
      WHEN  124 => Ti := "000001100100000110010001111110000010110010010111"; --    +410001    -512873
      WHEN  125 => Ti := "000001101111010100000100000010011101110111011100"; --    +455940    +646620
      WHEN  126 => Ti := "000010100111100011011001111101100101110001001000"; --    +686297    -631736
      WHEN  127 => Ti := "111010010001010101111001000001001001100110111101"; --   -1501831    +301501
      WHEN  128 => Ti := "000010010001010001110110000110000010011100001000"; --    +595062   +1582856
      WHEN  129 => Ti := "111100000111001001100010111101110110100001111010"; --   -1019294    -563078
      WHEN  130 => Ti := "111001010100011000011001111111110001100010110111"; --   -1751527     -59209
      WHEN  131 => Ti := "111110110010100111001000000000101001011010111110"; --    -316984    +169662
      WHEN  132 => Ti := "111110101010100101000010111011011000000010101101"; --    -349886   -1212243
      WHEN  133 => Ti := "000100101010100101110011111101110110110110110110"; --   +1223027    -561738
      WHEN  134 => Ti := "000101001111001110001010111000001000110010100000"; --   +1373066   -2061152
      WHEN  135 => Ti := "000000110000000100011101111111000111110001101100"; --    +196893    -230292
      WHEN  136 => Ti := "000010100101001101011111111100010001000110110000"; --    +676703    -978512
      WHEN  137 => Ti := "111110010011001100010011000001001011010111110010"; --    -445677    +308722
      WHEN  138 => Ti := "111100111100111010101110000000000010101010111001"; --    -799058     +10937
      WHEN  139 => Ti := "111111000111010110011110000000100011111011110110"; --    -232034    +147190
      WHEN  140 => Ti := "111100111000011101010001000001000010011000011100"; --    -817327    +271900
      WHEN  141 => Ti := "000011001000110111100001111101001111101111001000"; --    +822753    -721976
      WHEN  142 => Ti := "000100000010010111110101000011000000111101000001"; --   +1058293    +790337
      WHEN  143 => Ti := "111111111011000001001101000101000011101100000001"; --     -20403   +1325825
      WHEN  144 => Ti := "000000101000101010111011000011010111000100101111"; --    +166587    +880943
      WHEN  145 => Ti := "000000010101000110010010000100110000011011001111"; --     +86418   +1246927
      WHEN  146 => Ti := "111111001011110101011110000011110101011001111001"; --    -213666   +1005177
      WHEN  147 => Ti := "111001111001011110000011000001111011110001101111"; --   -1599613    +506991
      WHEN  148 => Ti := "000100010100010110111011111001101111010000000010"; --   +1131963   -1641470
      WHEN  149 => Ti := "111100111000000011111111111110011011011100101100"; --    -818945    -411860
      WHEN  150 => Ti := "111101011010000111101000000011011110100001001111"; --    -679448    +911439
      WHEN  151 => Ti := "000010110000000100010100111111001010000111010101"; --    +721172    -220715
      WHEN  152 => Ti := "000000101100001010110000000000011011101000101110"; --    +180912    +113198
      WHEN  153 => Ti := "000000100001000001111011111000011111010001001010"; --    +135291   -1969078
      WHEN  154 => Ti := "000001110010011001101110111101011001011000110001"; --    +468590    -682447
      WHEN  155 => Ti := "111110001011110000001101111110010011010010101110"; --    -476147    -445266
      WHEN  156 => Ti := "000000001110000111111000000100010010010100001000"; --     +57848   +1123592
      WHEN  157 => Ti := "000101000001111001000010000001010011100011010001"; --   +1318466    +342225
      WHEN  158 => Ti := "111100010110100001111000000011011100111011010001"; --    -956296    +904913
      WHEN  159 => Ti := "111110100111111000000010111110111001000011111011"; --    -360958    -290565
      WHEN  160 => Ti := "000011100011000111000110000001101010100110000100"; --    +930246    +436612
      WHEN  161 => Ti := "111111100111101100000010000100010001100111100000"; --     -99582   +1120736
      WHEN  162 => Ti := "111110100001000001011100111110100111011111110010"; --    -389028    -362510
      WHEN  163 => Ti := "111101100010100010011001000000111000100101011110"; --    -644967    +231774
      WHEN  164 => Ti := "111110000100111010010011111101101001101111010110"; --    -504173    -615466
      WHEN  165 => Ti := "000100001101111010001111000000110000111101111100"; --   +1105551    +200572
      WHEN  166 => Ti := "000000111011100011101001111100000100000101010011"; --    +243945   -1031853
      WHEN  167 => Ti := "000000011110011101100111000010001001010110101101"; --    +124775    +562605
      WHEN  168 => Ti := "000011000010011001011010000001110011001110100000"; --    +796250    +471968
      WHEN  169 => Ti := "000001111110001100001111000001011111110100011001"; --    +516879    +392473
      WHEN  170 => Ti := "111100101100100100100010000011001011101000000110"; --    -866014    +834054
      WHEN  171 => Ti := "000000010111001011011010000100001101100111011000"; --     +94938   +1104344
      WHEN  172 => Ti := "111101101000011110001011111010111111001100000110"; --    -620661   -1314042
      WHEN  173 => Ti := "000000011111011101110011000001000110110110100000"; --    +128883    +290208
      WHEN  174 => Ti := "000001001010000011010111111110011001110100110111"; --    +303319    -418505
      WHEN  175 => Ti := "000001010000000110001110111101011010001000101000"; --    +328078    -679384
      WHEN  176 => Ti := "000010111001011010110010000011001001011011010001"; --    +759474    +825041
      WHEN  177 => Ti := "111100101011000000001011000000001100011011110011"; --    -872437     +50931
      WHEN  178 => Ti := "111111110011101111110110000000111101010001000011"; --     -50186    +250947
      WHEN  179 => Ti := "000010101101101101011111111111101001111111111111"; --    +711519     -90113
      WHEN  180 => Ti := "000010000101101000000000000000001010000001111101"; --    +547328     +41085
      WHEN  181 => Ti := "111011111001111010001111000011100110110110001010"; --   -1073521    +945546
      WHEN  182 => Ti := "111110111000101001011110000001011111111101000110"; --    -292258    +393030
      WHEN  183 => Ti := "111110011011100000011101000001001111010011000011"; --    -411619    +324803
      WHEN  184 => Ti := "111100010011100010100101111100110000011011100011"; --    -968539    -850205
      WHEN  185 => Ti := "000000010110000101111110111100111101010001101111"; --     +90494    -797585
      WHEN  186 => Ti := "000000101100101111010010111110111101010000001100"; --    +183250    -273396
      WHEN  187 => Ti := "000000101000110110100001000000110110101001110100"; --    +167329    +223860
      WHEN  188 => Ti := "000000111010011010111001000001011000100011000101"; --    +239289    +362693
      WHEN  189 => Ti := "000011001100001100101111111110010110001010000011"; --    +836399    -433533
      WHEN  190 => Ti := "111100010011001111110010000010001110000010111001"; --    -969742    +581817
      WHEN  191 => Ti := "000011011001011101000011000010000011110000010010"; --    +890691    +539666
      WHEN  192 => Ti := "111100011000110001001010111011010100001010001001"; --    -947126   -1228151
      WHEN  193 => Ti := "111111111100101111011101000000100101000110110111"; --     -13347    +151991
      WHEN  194 => Ti := "111110010111111001110001000001001101000100010011"; --    -426383    +315667
      WHEN  195 => Ti := "000010001001011100100011000100000100100101101111"; --    +562979   +1067375
      WHEN  196 => Ti := "111110111101101100101110111111010111111000110001"; --    -271570    -164303
      WHEN  197 => Ti := "000010100011101010101110000000001101001010011110"; --    +670382     +53918
      WHEN  198 => Ti := "000010001011001001110100000000011010010000000011"; --    +569972    +107523
      WHEN  199 => Ti := "000101001011100001111000000000100110111010010000"; --   +1357944    +159376
      WHEN  200 => Ti := "111110000000110011001011111110001001101001111101"; --    -521013    -484739
      WHEN  201 => Ti := "111010000110010111001001111100110001001110001110"; --   -1546807    -846962
      WHEN  202 => Ti := "110100110110111111101001000010111010000111101111"; --   -2920471    +762351
      WHEN  203 => Ti := "111110101110010011010111111111100011001011010100"; --    -334633    -118060
      WHEN  204 => Ti := "111101010101001111110001111111110010001101001111"; --    -699407     -56497
      WHEN  205 => Ti := "111111111111101001001110000001000110111011100000"; --      -1458    +290528
      WHEN  206 => Ti := "000000000010000100101000000000111110100001010000"; --      +8488    +256080
      WHEN  207 => Ti := "000011111111010100001001000000001011000101010011"; --   +1045769     +45395
      WHEN  208 => Ti := "111101101000000100111001111101101111101110000010"; --    -622279    -590974
      WHEN  209 => Ti := "000001001000000100100011000010000101110110000100"; --    +295203    +548228
      WHEN  210 => Ti := "111111111101111000110001111111001000010000011010"; --      -8655    -228326
      WHEN  211 => Ti := "000000001010011110100111111110000001000111001111"; --     +42919    -519729
      WHEN  212 => Ti := "000000110101001001100001000010110010110001011010"; --    +217697    +732250
      WHEN  213 => Ti := "110111011010011001000011111110110101110110111110"; --   -2251197    -303682
      WHEN  214 => Ti := "111111001000000001100000111101011111100111101000"; --    -229280    -656920
      WHEN  215 => Ti := "000100110110101101010110111110001000100011010101"; --   +1272662    -489259
      WHEN  216 => Ti := "000101011010101100000001000011011110011101000110"; --   +1420033    +911174
      WHEN  217 => Ti := "111110101100100100101111000001100000010011011011"; --    -341713    +394459
      WHEN  218 => Ti := "111101110111111000010001111100110011000110011000"; --    -557551    -839272
      WHEN  219 => Ti := "000110110001111111101011000010010001111011010111"; --   +1777643    +597719
      WHEN  220 => Ti := "000001000100101111000111000101001011001001010110"; --    +281543   +1356374
      WHEN  221 => Ti := "111111110111000000111001111011010100110110101000"; --     -36807   -1225304
      WHEN  222 => Ti := "111100111110110100111101000000110110111101101100"; --    -791235    +225132
      WHEN  223 => Ti := "000001001111110101011101111111100000001110010001"; --    +327005    -130159
      WHEN  224 => Ti := "000011100010001000011101000010111000111101111110"; --    +926237    +757630
      WHEN  225 => Ti := "111101011001101001110010111111111101001101000100"; --    -681358     -11452
      WHEN  226 => Ti := "000001010000011101100100111011110001101111000100"; --    +329572   -1107004
      WHEN  227 => Ti := "000000010010000000100101000001001001000111101111"; --     +73765    +299503
      WHEN  228 => Ti := "000001100110111011011101111101101110100110001010"; --    +421597    -595574
      WHEN  229 => Ti := "111010111010101101011001111110100110010001010010"; --   -1332391    -367534
      WHEN  230 => Ti := "111011100010011011111111111011011010000110110001"; --   -1169665   -1203791
      WHEN  231 => Ti := "000011101111100010111001111101000010010001010010"; --    +981177    -777134
      WHEN  232 => Ti := "000000010000000110101010111100010111100001010011"; --     +65962    -952237
      WHEN  233 => Ti := "000001100010111111110010111111001011000101001111"; --    +405490    -216753
      WHEN  234 => Ti := "111111100011000101011101000000011110101100011001"; --    -118435    +125721
      WHEN  235 => Ti := "111110000110000010111100111110101111101111011010"; --    -499524    -328742
      WHEN  236 => Ti := "000000100111100110100000000001010001011000001000"; --    +162208    +333320
      WHEN  237 => Ti := "111111010110010001010100111110100111001011010010"; --    -170924    -363822
      WHEN  238 => Ti := "111011101110011111001011000000010001111111100010"; --   -1120309     +73698
      WHEN  239 => Ti := "111111110101000100001001111010001000011100101111"; --     -44791   -1538257
      WHEN  240 => Ti := "111110100101111010010011111110011110101100110010"; --    -369005    -398542
      WHEN  241 => Ti := "000011010011101001011110000001110011001010011011"; --    +866910    +471707
      WHEN  242 => Ti := "000000111000000000101110111111101100001100001111"; --    +229422     -81137
      WHEN  243 => Ti := "111110011110000101100000111111011101111111101000"; --    -401056    -139288
      WHEN  244 => Ti := "111111101011010111011011111111110010001001001110"; --     -84517     -56754
      WHEN  245 => Ti := "111110010001000100000101000001111000000111110000"; --    -454395    +492016
      WHEN  246 => Ti := "000010111111100111001111000011000010100111101101"; --    +784847    +797165
      WHEN  247 => Ti := "111001011010011111110111111111011010000011101000"; --   -1726473    -155416
      WHEN  248 => Ti := "111110000010000011001111111110011010010100111110"; --    -515889    -416450
      WHEN  249 => Ti := "111111100101110000011001000010011011010111100011"; --    -107495    +636387
      WHEN  250 => Ti := "111111011011011001111111000001111101010000010011"; --    -149889    +513043
      WHEN  251 => Ti := "111110011101110000101101111100000011111010001110"; --    -402387   -1032562
      WHEN  252 => Ti := "000101110101011111001011111110101101111010011111"; --   +1529803    -336225
      WHEN  253 => Ti := "111111100011010000001100000101011001001111110101"; --    -117748   +1414133
      WHEN  254 => Ti := "000000100010010011001100000000100001101100101000"; --    +140492    +138024
      WHEN  255 => Ti := "111100010010111010011101000000010000100011010010"; --    -971107     +67794
      WHEN  256 => Ti := "000100101000100000001100111111000000011010101001"; --   +1214476    -260439
      WHEN  257 => Ti := "000000101110100001110000111101101000111111001110"; --    +190576    -618546
      WHEN  258 => Ti := "111100110100110000110100111010111011110101001111"; --    -832460   -1327793
      WHEN  259 => Ti := "000010000001100000101000111101110110100011110101"; --    +530472    -562955
      WHEN  260 => Ti := "111101110101100100111010111111110111011011000111"; --    -566982     -35129
      WHEN  261 => Ti := "111101010010001010001000111110110001010111110100"; --    -712056    -322060
      WHEN  262 => Ti := "111101111101010110011001111101000010111010111111"; --    -535143    -774465
      WHEN  263 => Ti := "111100010001001111110101000010101110001010101011"; --    -977931    +713387
      WHEN  264 => Ti := "111110110011010001100110111110111100010011001011"; --    -314266    -277301
      WHEN  265 => Ti := "000000110110010100000000000000010001000010111011"; --    +222464     +69819
      WHEN  266 => Ti := "111110010000001001110100111011011011101101110000"; --    -458124   -1197200
      WHEN  267 => Ti := "111110000010000111001110111101010110011100001001"; --    -515634    -694519
      WHEN  268 => Ti := "000001110011101011001011111110110001111000011011"; --    +473803    -319973
      WHEN  269 => Ti := "111011000000001100111110000000000001110011000010"; --   -1309890      +7362
      WHEN  270 => Ti := "000000111010001111111011111110000000001010111110"; --    +238587    -523586
      WHEN  271 => Ti := "111110100000110011000111111101100001011011110100"; --    -389945    -649484
      WHEN  272 => Ti := "111100110101101001010111000101100101001101100111"; --    -828841   +1463143
      WHEN  273 => Ti := "111110111011000001010000000000111011111100010001"; --    -282544    +245521
      WHEN  274 => Ti := "111011101100000111111100000010111010101010010001"; --   -1129988    +764561
      WHEN  275 => Ti := "000000111010010011000001111100100100111011110101"; --    +238785    -897291
      WHEN  276 => Ti := "000001100111011101110101000001100110011101110101"; --    +423797    +419701
      WHEN  277 => Ti := "111111100011001010011100000000011001100000111010"; --    -118116    +104506
      WHEN  278 => Ti := "111010101001001110010101000011110000110000000010"; --   -1404011    +986114
      WHEN  279 => Ti := "111101101011111000010100000010100101010110111010"; --    -606700    +677306
      WHEN  280 => Ti := "111110100110011011010101000101111110010101110001"; --    -366891   +1566065
      WHEN  281 => Ti := "111110011110000100011110111110100101000100010000"; --    -401122    -372464
      WHEN  282 => Ti := "000000001110100010001100111111101010011001000001"; --     +59532     -88511
      WHEN  283 => Ti := "000000111111011110000100000000110101011101100010"; --    +259972    +218978
      WHEN  284 => Ti := "000100100010000101000010111111111010011111100001"; --   +1188162     -22559
      WHEN  285 => Ti := "111100110100001100010111111110110101001000010111"; --    -834793    -306665
      WHEN  286 => Ti := "111110101000001101111001111111111011101000111110"; --    -359559     -17858
      WHEN  287 => Ti := "111111011101001100010101111011001100100100110000"; --    -142571   -1259216
      WHEN  288 => Ti := "111111100101110111010101000001100111111111101010"; --    -107051    +425962
      WHEN  289 => Ti := "000001001110111101100010111110010111110011100100"; --    +323426    -426780
      WHEN  290 => Ti := "000010000111100011001101111011001111010010001100"; --    +555213   -1248116
      WHEN  291 => Ti := "000001011011100001110110111011011100110100001011"; --    +374902   -1192693
      WHEN  292 => Ti := "111101001010111011100011000000011110001111101000"; --    -741661    +123880
      WHEN  293 => Ti := "111101110101000111101110000010000110111010110000"; --    -568850    +552624
      WHEN  294 => Ti := "000100011101011000101101000010101111111011000111"; --   +1168941    +720583
      WHEN  295 => Ti := "000001111010011100000110111111010110101110011010"; --    +501510    -169062
      WHEN  296 => Ti := "111111010101011110011011000000100101001001000000"; --    -174181    +152128
      WHEN  297 => Ti := "000110111111001100111100000010100010000100000101"; --   +1831740    +663813
      WHEN  298 => Ti := "000000010011110100000101000000010110111010101111"; --     +81157     +93871
      WHEN  299 => Ti := "000100100011110010010000000000000011110100010100"; --   +1195152     +15636
      WHEN  300 => Ti := "000001001010000100110100111110010100111001010010"; --    +303412    -438702
      WHEN  301 => Ti := "111011100000111100100011111011000101101000000011"; --   -1175773   -1287677
      WHEN  302 => Ti := "000000111000000000110010111111100101110111010110"; --    +229426    -107050
      WHEN  303 => Ti := "000000001110000011110101111110100000001111011101"; --     +57589    -392227
      WHEN  304 => Ti := "111110110000101010010100111111101110000001111100"; --    -324972     -73604
      WHEN  305 => Ti := "111101100101101111111110000000000111001010000110"; --    -631810     +29318
      WHEN  306 => Ti := "111101001000011110001000000100111100100011101001"; --    -751736   +1296617
      WHEN  307 => Ti := "111101100011100101010010111011111000011101100011"; --    -640686   -1079453
      WHEN  308 => Ti := "000010110111110110010111000000010111011010110111"; --    +753047     +95927
      WHEN  309 => Ti := "111110001110110110111110000010000010110010011001"; --    -463426    +535705
      WHEN  310 => Ti := "111110110011111101001001111110011110111001001111"; --    -311479    -397745
      WHEN  311 => Ti := "000011111100010111011110111111111111011101010001"; --   +1033694      -2223
      WHEN  312 => Ti := "000010111111100010011100000011010101011011110110"; --    +784540    +874230
      WHEN  313 => Ti := "111111011101110001011001111100101101101110001100"; --    -140199    -861300
      WHEN  314 => Ti := "000000100111010100001111000001000010111110000001"; --    +161039    +274305
      WHEN  315 => Ti := "111110111000011000111011111111100111000001101001"; --    -293317    -102295
      WHEN  316 => Ti := "111010110001011000010100111110100100010001100010"; --   -1370604    -375710
      WHEN  317 => Ti := "000011011000110100000100000010100000001010000000"; --    +888068    +656000
      WHEN  318 => Ti := "111110011001010111001001111000100111101101011011"; --    -420407   -1934501
      WHEN  319 => Ti := "000000001001111010111000111100001011001110000011"; --     +40632   -1002621
      WHEN  320 => Ti := "000000011111000001000101000001010010100000000111"; --    +127045    +337927
      WHEN  321 => Ti := "111111101010111111010101111101101110001000111110"; --     -86059    -597442
      WHEN  322 => Ti := "111111100100101001111111000010000101101101000100"; --    -112001    +547652
      WHEN  323 => Ti := "000000000100111100000010000001000100011001001111"; --     +20226    +280143
      WHEN  324 => Ti := "111111110001110111101110111011111011101111011101"; --     -57874   -1066019
      WHEN  325 => Ti := "111111010101100100110010111110001111111111100110"; --    -173774    -458778
      WHEN  326 => Ti := "111100110110011101010011111111001000111011011011"; --    -825517    -225573
      WHEN  327 => Ti := "000001000010111010000111000110110011010000011111"; --    +274055   +1782815
      WHEN  328 => Ti := "111101111000011001111100000011100101010100000011"; --    -555396    +939267
      WHEN  329 => Ti := "000000110111100001111010000000101010010110100100"; --    +227450    +173476
      WHEN  330 => Ti := "111111000001111100010110000010011010010000010111"; --    -254186    +631831
      WHEN  331 => Ti := "000010011110110011111101000011010110000110010111"; --    +650493    +876951
      WHEN  332 => Ti := "000000111001110100110010000001011000100000100000"; --    +236850    +362528
      WHEN  333 => Ti := "000000011101100001100110000000100111111001010000"; --    +120934    +163408
      WHEN  334 => Ti := "111100101111010110000000111111000000001100000100"; --    -854656    -261372
      WHEN  335 => Ti := "111100100000111000101101111111110011101111111000"; --    -913875     -50184
      WHEN  336 => Ti := "111111111010111101000011000000100101010011111010"; --     -20669    +152826
      WHEN  337 => Ti := "111111100100111111001000000010111000000010110000"; --    -110648    +753840
      WHEN  338 => Ti := "111111100011100001101110000111010110011100011110"; --    -116626   +1926942
      WHEN  339 => Ti := "111111001101111000000000000010011100110010010010"; --    -205312    +642194
      WHEN  340 => Ti := "000011101110110000011001000011010110010000101011"; --    +977945    +877611
      WHEN  341 => Ti := "000001100111001000011101000101100110010110011110"; --    +422429   +1467806
      WHEN  342 => Ti := "000100011110011110110101111101001010110111100111"; --   +1173429    -741913
      WHEN  343 => Ti := "111011001110001010110011111110011011011001101001"; --   -1252685    -412055
      WHEN  344 => Ti := "000001101011000001101101000001010111110010101010"; --    +438381    +359594
      WHEN  345 => Ti := "000010001001110101011110111100010011011110000110"; --    +564574    -968826
      WHEN  346 => Ti := "111111010101001010111000000000000101111100001000"; --    -175432     +24328
      WHEN  347 => Ti := "000001111001111100010111000011011000011101001010"; --    +499479    +886602
      WHEN  348 => Ti := "111110101000100001110100000010111001111001100101"; --    -358284    +761445
      WHEN  349 => Ti := "000000110111010101011101111001111100111010011110"; --    +226653   -1585506
      WHEN  350 => Ti := "111111101110100001000110111110111101100011011100"; --     -71610    -272164
      WHEN  351 => Ti := "111101101010101010001110111011101011011100011010"; --    -611698   -1132774
      WHEN  352 => Ti := "111101110100110100010100111101101001111000000000"; --    -570092    -614912
      WHEN  353 => Ti := "111100010100110011101001000010111100001001001011"; --    -963351    +770635
      WHEN  354 => Ti := "111100100011010101101001000001011001101101111000"; --    -903831    +367480
      WHEN  355 => Ti := "111101111001000110111011000010001100001101010001"; --    -552517    +574289
      WHEN  356 => Ti := "000010110101001110001100111101011000101000011001"; --    +742284    -685543
      WHEN  357 => Ti := "111010101111011000000001000010000011111111011100"; --   -1378815    +540636
      WHEN  358 => Ti := "111111100111101011110011111110110101011110001001"; --     -99597    -305271
      WHEN  359 => Ti := "111111101000100100101010000000101101010110100100"; --     -95958    +185764
      WHEN  360 => Ti := "000010100100010110001010111101000001111100100001"; --    +673162    -778463
      WHEN  361 => Ti := "111111011101000000111011111100111001001101110010"; --    -143301    -814222
      WHEN  362 => Ti := "111100000001100101111011111110101101011010110001"; --   -1042053    -338255
      WHEN  363 => Ti := "111111100010101011001111111100001110111101010001"; --    -120113    -987311
      WHEN  364 => Ti := "000010001110100000000011111111011111011001100101"; --    +583683    -133531
      WHEN  365 => Ti := "000011101001101001000000000001000001001111011101"; --    +956992    +267229
      WHEN  366 => Ti := "111110110110000100111001111110110010100010010111"; --    -302791    -317289
      WHEN  367 => Ti := "000100001100101111100000000001100000011110001100"; --   +1100768    +395148
      WHEN  368 => Ti := "111111010111001001011100000001010110010010000001"; --    -167332    +353409
      WHEN  369 => Ti := "000000000111100000001011111100111111010000001101"; --     +30731    -789491
      WHEN  370 => Ti := "000001100110010010001101000001110001010100111110"; --    +418957    +464190
      WHEN  371 => Ti := "000010111110010111111101000010111000010011010111"; --    +779773    +754903
      WHEN  372 => Ti := "111111110110111010001011111110011000101101101011"; --     -37237    -423061
      WHEN  373 => Ti := "000001000011000010110101000001101111111000110011"; --    +274613    +458291
      WHEN  374 => Ti := "000000111010101001100000111110111010101010001111"; --    +240224    -284017
      WHEN  375 => Ti := "000001101111000100111110000000101011110110011000"; --    +454974    +179608
      WHEN  376 => Ti := "000000111111111101001110111110001110111100000111"; --    +261966    -463097
      WHEN  377 => Ti := "111111110101010001111100111100011010111100000110"; --     -43908    -938234
      WHEN  378 => Ti := "000010010110100111000111111100111110001011100010"; --    +616903    -793886
      WHEN  379 => Ti := "000101101111000110100110111101000001010000100101"; --   +1503654    -781275
      WHEN  380 => Ti := "000001000111111001010010000000111100100111010010"; --    +294482    +248274
      WHEN  381 => Ti := "111111111010011101010000111100100001100111100110"; --     -22704    -910874
      WHEN  382 => Ti := "000010101101010110010001111110101010100101101110"; --    +710033    -349842
      WHEN  383 => Ti := "111110100110001110000101000001011111010000100001"; --    -367739    +390177
      WHEN  384 => Ti := "000000001100110010011111111010100010000110101001"; --     +52383   -1433175
      WHEN  385 => Ti := "111011011001011011111010111110110101111100111110"; --   -1206534    -303298
      WHEN  386 => Ti := "111101011011111111101010111010101000111110011011"; --    -671766   -1405029
      WHEN  387 => Ti := "000010100000110000100101111111101010111010110000"; --    +658469     -86352
      WHEN  388 => Ti := "111110111100010101110110111111010000001100110101"; --    -277130    -195787
      WHEN  389 => Ti := "000001011111100010000000000010101011011111100011"; --    +391296    +702435
      WHEN  390 => Ti := "000000110100001100101101111111100001000110100101"; --    +213805    -126555
      WHEN  391 => Ti := "111110010101000111010001111110001101010100101010"; --    -437807    -469718
      WHEN  392 => Ti := "000010010011001111111100111101000011111111100010"; --    +603132    -770078
      WHEN  393 => Ti := "111100001111101100000000111101101110001011111010"; --    -984320    -597254
      WHEN  394 => Ti := "111101001111101011100010111100100001001111010001"; --    -722206    -912431
      WHEN  395 => Ti := "000001001000111100000001000101110010011111101100"; --    +298753   +1517548
      WHEN  396 => Ti := "000011001011110110010001111110111011000110001101"; --    +834961    -282227
      WHEN  397 => Ti := "111111110110001011101111000011011011100111101010"; --     -40209    +899562
      WHEN  398 => Ti := "000001101100010111100001000100001010111000111010"; --    +443873   +1093178
      WHEN  399 => Ti := "111111011111111110100001111110100011001100001101"; --    -131167    -380147
      WHEN  400 => Ti := "000000100111011010011100000000011001111011111011"; --    +161436    +106235
      WHEN  401 => Ti := "111110100100000101011011111111001101110100010111"; --    -376485    -205545
      WHEN  402 => Ti := "000001100000011110110101111111100001001101011110"; --    +395189    -126114
      WHEN  403 => Ti := "000000111001000101100110111111001010100011001000"; --    +233830    -218936
      WHEN  404 => Ti := "000011010101010101010110111110100100110111011000"; --    +873814    -373288
      WHEN  405 => Ti := "000001100101110110110100111011100000010000001001"; --    +417204   -1178615
      WHEN  406 => Ti := "000001011001010100011000000000101001100010110001"; --    +365848    +170161
      WHEN  407 => Ti := "000010010010000001100010000001101110100001101000"; --    +598114    +452712
      WHEN  408 => Ti := "000000001011010110101111000000011001000010010001"; --     +46511    +102545
      WHEN  409 => Ti := "111101000100000001110111000000010111110100111100"; --    -769929     +97596
      WHEN  410 => Ti := "111101101010101101111001000000010100100001001110"; --    -611463     +84046
      WHEN  411 => Ti := "111101011111101111010011000101100000111101000100"; --    -656429   +1445700
      WHEN  412 => Ti := "111111101111100111110110111101000111000100101011"; --     -67082    -757461
      WHEN  413 => Ti := "000001000110100010010010111111101100010011010101"; --    +288914     -80683
      WHEN  414 => Ti := "111010101001000011110111111101110011001110010100"; --   -1404681    -576620
      WHEN  415 => Ti := "111111101100110111100000000010010101000000011101"; --     -78368    +610333
      WHEN  416 => Ti := "111111110111111100111001000011010010000011111011"; --     -32967    +860411
      WHEN  417 => Ti := "111111110010101011010000111111001100010111001010"; --     -54576    -211510
      WHEN  418 => Ti := "111111100110111001010000111110100110000010000011"; --    -102832    -368509
      WHEN  419 => Ti := "111110000110010000011110000010011010111011111110"; --    -498658    +634622
      WHEN  420 => Ti := "111111101001010100001100000001110101111101100111"; --     -92916    +483175
      WHEN  421 => Ti := "000000101011010111111010000000111110100100101011"; --    +177658    +256299
      WHEN  422 => Ti := "111111110001110000110001000111011011110000100111"; --     -58319   +1948711
      WHEN  423 => Ti := "000000100011001101110010000001001110100110000100"; --    +144242    +321924
      WHEN  424 => Ti := "000100010001011001110001000001000101001110001111"; --   +1119857    +283535
      WHEN  425 => Ti := "111010001101001000011110000101000110110101101111"; --   -1519074   +1338735
      WHEN  426 => Ti := "000001001110001110110010000100010111111110010001"; --    +320434   +1146769
      WHEN  427 => Ti := "111100110000110101111101111101110000010010011010"; --    -848515    -588646
      WHEN  428 => Ti := "111100110100000011001001000100110000001111101100"; --    -835383   +1246188
      WHEN  429 => Ti := "111101110100000101100100111110100100010110110101"; --    -573084    -375371
      WHEN  430 => Ti := "111110110000010000010100111110001100110000001000"; --    -326636    -472056
      WHEN  431 => Ti := "111110110000001010010110111110100011100000000110"; --    -327018    -378874
      WHEN  432 => Ti := "000001100011111011011010000000001011011110100110"; --    +409306     +47014
      WHEN  433 => Ti := "000100000111011011100000111100111111000000000110"; --   +1079008    -790522
      WHEN  434 => Ti := "000001100111111000000010111111110011001010100111"; --    +425474     -52569
      WHEN  435 => Ti := "111011111100010111011011111011100111101100100011"; --   -1063461   -1148125
      WHEN  436 => Ti := "111101011100110100011001000100000111111000101011"; --    -668391   +1080875
      WHEN  437 => Ti := "111110111110110001110101111011111000110111111001"; --    -267147   -1077767
      WHEN  438 => Ti := "000000110000110101110010111101100110011111001010"; --    +200050    -628790
      WHEN  439 => Ti := "111101111110011011011001000000100110100010010101"; --    -530727    +157845
      WHEN  440 => Ti := "000000100000000010101001111110001001001100111101"; --    +131241    -486595
      WHEN  441 => Ti := "111111010110011111100000000000010011010111010000"; --    -170016     +79312
      WHEN  442 => Ti := "111111010000001111110000000001000000001011000101"; --    -195600    +262853
      WHEN  443 => Ti := "111010101101101100000110111110100000111011111011"; --   -1385722    -389381
      WHEN  444 => Ti := "000000100101011011001011000010011001101010101010"; --    +153291    +629418
      WHEN  445 => Ti := "000010010001000010100001111111101001000100011110"; --    +594081     -93922
      WHEN  446 => Ti := "111110110110100111011110111111011101011001101011"; --    -300578    -141717
      WHEN  447 => Ti := "000001110001011010101100000010110111001001010000"; --    +464556    +750160
      WHEN  448 => Ti := "111111011010000100001010111100110100010110000001"; --    -155382    -834175
      WHEN  449 => Ti := "000000010110111001000101000001001011001011011110"; --     +93765    +307934
      WHEN  450 => Ti := "000011100000110000101111111111111111010111001001"; --    +920623      -2615
      WHEN  451 => Ti := "111111100011000000111111000001000100101110110110"; --    -118721    +281526
      WHEN  452 => Ti := "000001100110011110101010111101001101110001110011"; --    +419754    -729997
      WHEN  453 => Ti := "111101010100111000001111000000101011101000001111"; --    -700913    +178703
      WHEN  454 => Ti := "000000010111001010000011000110100001001011011001"; --     +94851   +1708761
      WHEN  455 => Ti := "000001000110001101111000000000100001011011001000"; --    +287608    +136904
      WHEN  456 => Ti := "000001111100101000100111000000101011011101111000"; --    +510503    +178040
      WHEN  457 => Ti := "000001100100101110100111111101011011001000110110"; --    +412583    -675274
      WHEN  458 => Ti := "000000001110110010011011000001110110100101111110"; --     +60571    +485758
      WHEN  459 => Ti := "000000110111010110001110000000001010010011001000"; --    +226702     +42184
      WHEN  460 => Ti := "111100100001111110010010000000111011000001000111"; --    -909422    +241735
      WHEN  461 => Ti := "000010001001000001110110000010101101110000001011"; --    +561270    +711691
      WHEN  462 => Ti := "000010010011101100001001000011100100000010001001"; --    +604937    +934025
      WHEN  463 => Ti := "000000101111011010001000111110111011110010010011"; --    +194184    -279405
      WHEN  464 => Ti := "111111000101111011100111000100011100010011001011"; --    -237849   +1164491
      WHEN  465 => Ti := "000000110001101000010011000000101000110111010101"; --    +203283    +167381
      WHEN  466 => Ti := "000000101110000010011001111101000101001101001011"; --    +188569    -765109
      WHEN  467 => Ti := "111111101100111000100111000001001000011010010111"; --     -78297    +296599
      WHEN  468 => Ti := "000000000111010001111111000001010111110010110000"; --     +29823    +359600
      WHEN  469 => Ti := "111110100111101001101000111111000010010011101011"; --    -361880    -252693
      WHEN  470 => Ti := "111111110001111010111011000010001001111011001101"; --     -57669    +564941
      WHEN  471 => Ti := "000000000001000011011101111110110001011001011001"; --      +4317    -321959
      WHEN  472 => Ti := "000001000101011111001000111111000100001011111110"; --    +284616    -244994
      WHEN  473 => Ti := "111111111100111111001110111110110100000010101110"; --     -12338    -311122
      WHEN  474 => Ti := "111111000100011111001110111100000110010001101110"; --    -243762   -1022866
      WHEN  475 => Ti := "111101101110110001100110000001101010000101010110"; --    -594842    +434518
      WHEN  476 => Ti := "000000000011000110101010111001111000111010100010"; --     +12714   -1601886
      WHEN  477 => Ti := "000000011000101011110001111011110010011010110001"; --    +101105   -1104207
      WHEN  478 => Ti := "000011110100010111010110111111100001100010011111"; --   +1000918    -124769
      WHEN  479 => Ti := "111101110110100100101011000010100000010110101001"; --    -562901    +656809
      WHEN  480 => Ti := "111110011010111101011001000001010101011010110101"; --    -413863    +349877
      WHEN  481 => Ti := "000000110011001011111011000001111111001111001111"; --    +209659    +521167
      WHEN  482 => Ti := "000011101011111011110000000110001010101101011111"; --    +966384   +1616735
      WHEN  483 => Ti := "111110011110011001010111111111100111111100011001"; --    -399785     -98535
      WHEN  484 => Ti := "111110111010110110011001111001111011000000101101"; --    -283239   -1593299
      WHEN  485 => Ti := "000011000001010100110100111111110001011100001111"; --    +791860     -59633
      WHEN  486 => Ti := "111100100000010100100011000011001001111011101101"; --    -916189    +827117
      WHEN  487 => Ti := "000010000011001001110010111101111000111010100110"; --    +537202    -553306
      WHEN  488 => Ti := "000011000000010010111100111110001000001010011001"; --    +787644    -490855
      WHEN  489 => Ti := "000011001100000110001111000001100100011101000000"; --    +835983    +411456
      WHEN  490 => Ti := "111110001011001011000011111011101010000011101110"; --    -478525   -1138450
      WHEN  491 => Ti := "111011101100001110001111000000011110000010010001"; --   -1129585    +123025
      WHEN  492 => Ti := "111110100011001110011101000000000101010100010100"; --    -380003     +21780
      WHEN  493 => Ti := "111111100010100111010011111101111101110010100010"; --    -120365    -533342
      WHEN  494 => Ti := "000011100110101110011001111111100111101011111110"; --    +945049     -99586
      WHEN  495 => Ti := "111111101111100100011000000001111000000000101110"; --     -67304    +491566
      WHEN  496 => Ti := "111011100110100000111010000001110001101101100001"; --   -1152966    +465761
      WHEN  497 => Ti := "111100110010000001010111000101011010110101100100"; --    -843689   +1420644
      WHEN  498 => Ti := "000011011011010111101111000011100000000010000001"; --    +898543    +917633
      WHEN  499 => Ti := "111100101100111111101000000100100100011101001101"; --    -864280   +1197901
      WHEN  500 => Ti := "000000011101001110100110111111101010110111111110"; --    +119718     -86530
      WHEN  501 => Ti := "000010100100011001110111000000111111000010010101"; --    +673399    +258197
      WHEN  502 => Ti := "000011111000100101101111000001011101000101010110"; --   +1018223    +381270
      WHEN  503 => Ti := "111110010101101101010110000000000100100100001011"; --    -435370     +18699
      WHEN  504 => Ti := "111001100011101001000110000001101010110111010100"; --   -1689018    +437716
      WHEN  505 => Ti := "000011100000010111100011000000000010100110110011"; --    +919011     +10675
      WHEN  506 => Ti := "000000100000011111001100000000011110110011101010"; --    +133068    +126186
      WHEN  507 => Ti := "111011000111010101011111111100000010100000001101"; --   -1280673   -1038323
      WHEN  508 => Ti := "000001010100011001001100111111010111110011000000"; --    +345676    -164672
      WHEN  509 => Ti := "000001111000011000101011000001110001000011001000"; --    +493099    +463048
      WHEN  510 => Ti := "111011111000010010101001111111010011110000000100"; --   -1080151    -181244
      WHEN  511 => Ti := "000001000111001110101000000100010101001000010100"; --    +291752   +1135124
      WHEN  512 => Ti := "111111000000100101000111111111111111010111101000"; --    -259769      -2584
      WHEN  513 => Ti := "111011011101110000100000000100010100100101100100"; --   -1188832   +1132900
      WHEN  514 => Ti := "111111101001111010011100111110000101110110010011"; --     -90468    -500333
      WHEN  515 => Ti := "111110111010111010010101111110011000000101010110"; --    -282987    -425642
      WHEN  516 => Ti := "000000011110001111100001000000010110110011001100"; --    +123873     +93388
      WHEN  517 => Ti := "111111010101000101101111000010011101100001011001"; --    -175761    +645209
      WHEN  518 => Ti := "000001110010110111100011000011111110010100011010"; --    +470499   +1041690
      WHEN  519 => Ti := "000001111001010110000000000000000011010011100011"; --    +497024     +13539
      WHEN  520 => Ti := "111110001000000011111100000001000111101101111111"; --    -491268    +293759
      WHEN  521 => Ti := "111100110110111000110000111111101010111111111111"; --    -823760     -86017
      WHEN  522 => Ti := "000001001101001100001010111011100110011101000101"; --    +316170   -1153211
      WHEN  523 => Ti := "000011001011101111010000111100111111010100101111"; --    +834512    -789201
      WHEN  524 => Ti := "111111010100111101110110111111001011010010010111"; --    -176266    -215913
      WHEN  525 => Ti := "000000110001011010010011000000111010011000000011"; --    +202387    +239107
      WHEN  526 => Ti := "000000010011110110011010111110110100000100111000"; --     +81306    -310984
      WHEN  527 => Ti := "111110010100001000110001111111010011111100111111"; --    -441807    -180417
      WHEN  528 => Ti := "111110111010010111000110111101100000001010010001"; --    -285242    -654703
      WHEN  529 => Ti := "111110010001000100000110111110101010100100110011"; --    -454394    -349901
      WHEN  530 => Ti := "000001111100101110010100000011000111000111101101"; --    +510868    +815597
      WHEN  531 => Ti := "000010111111101001000000111111111001101110000110"; --    +784960     -25722
      WHEN  532 => Ti := "111111000010010101101100111101001110000000101011"; --    -252564    -729045
      WHEN  533 => Ti := "000011010011010000010100000000111100111111111100"; --    +865300    +249852
      WHEN  534 => Ti := "000101001101000001111110000010111111101011101010"; --   +1364094    +785130
      WHEN  535 => Ti := "000111001010110011011011000101100010001000101110"; --   +1879259   +1450542
      WHEN  536 => Ti := "111110100001010100111100000011011100110110010011"; --    -387780    +904595
      WHEN  537 => Ti := "111100111100010000111011000011000000000111000100"; --    -801733    +786884
      WHEN  538 => Ti := "111111001100000000100000111111100000101000001110"; --    -212960    -128498
      WHEN  539 => Ti := "111111100110100010110100000001010111010100011000"; --    -104268    +357656
      WHEN  540 => Ti := "000000010000011010110000111101010111001111011110"; --     +67248    -691234
      WHEN  541 => Ti := "111111110000010000111010000000100001101111000010"; --     -64454    +138178
      WHEN  542 => Ti := "000000001111111001011111000001110010000110101111"; --     +65119    +467375
      WHEN  543 => Ti := "111100001000100000001101000010110110101011001011"; --   -1013747    +748235
      WHEN  544 => Ti := "000001000111101000010110111101010100111011000000"; --    +293398    -700736
      WHEN  545 => Ti := "000010000000110000101000111100011011001100010001"; --    +527400    -937199
      WHEN  546 => Ti := "111111101110000110011100111010010000111100111010"; --     -73316   -1503430
      WHEN  547 => Ti := "111111101110110001111000000001101001001010000010"; --     -70536    +430722
      WHEN  548 => Ti := "111000111100111111010011000100011100010011111110"; --   -1847341   +1164542
      WHEN  549 => Ti := "000011010110110001010000111100100000110110101010"; --    +879696    -914006
      WHEN  550 => Ti := "000000100101111001000110000000010011100101100011"; --    +155206     +80227
      WHEN  551 => Ti := "111111000010110010110100000000100101001001001111"; --    -250700    +152143
      WHEN  552 => Ti := "111110111100010110111001111110111111110111010001"; --    -277063    -262703
      WHEN  553 => Ti := "000010000011101000011111111110111001001000001100"; --    +539167    -290292
      WHEN  554 => Ti := "111110010011110101010000000001000100110011110000"; --    -443056    +281840
      WHEN  555 => Ti := "000000001000100101010000000001110110011010011100"; --     +35152    +485020
      WHEN  556 => Ti := "000011100000111111011110111111001011100010011111"; --    +921566    -214881
      WHEN  557 => Ti := "000110001001010110110111000011100110010010111110"; --   +1611191    +943294
      WHEN  558 => Ti := "111110001001100110001100000010001100010001000110"; --    -484980    +574534
      WHEN  559 => Ti := "000101100111110100011000111111100011111110110001"; --   +1473816    -114767
      WHEN  560 => Ti := "000011100011110100100101000110010100001110001000"; --    +933157   +1655688
      WHEN  561 => Ti := "000010111101111010000011000001000010100011110010"; --    +777859    +272626
      WHEN  562 => Ti := "111111010100100011010001111100111010100110010111"; --    -177967    -808553
      WHEN  563 => Ti := "000010100100011000111001000001000001000100111000"; --    +673337    +266552
      WHEN  564 => Ti := "111110011101001001110100111111010101011011110010"; --    -404876    -174350
      WHEN  565 => Ti := "111101101010011010101010000000011100010011010000"; --    -612694    +115920
      WHEN  566 => Ti := "111100001001010101010000000010111000100100100000"; --   -1010352    +756000
      WHEN  567 => Ti := "000000110101010100111011111010011100110111101111"; --    +218427   -1454609
      WHEN  568 => Ti := "111110011111111110110111000001001111101001000101"; --    -393289    +326213
      WHEN  569 => Ti := "000010110000011011100010111111011011100000111001"; --    +722658    -149447
      WHEN  570 => Ti := "000001011001001110011101111111100011000110001111"; --    +365469    -118385
      WHEN  571 => Ti := "111110101001101010011001111111111001010111100010"; --    -353639     -27166
      WHEN  572 => Ti := "000101001111011001111101111110110100100000110011"; --   +1373821    -309197
      WHEN  573 => Ti := "000010011100011000001011111111011000111111101111"; --    +640523    -159761
      WHEN  574 => Ti := "000101111100001101001111111101011010101101011010"; --   +1557327    -677030
      WHEN  575 => Ti := "000001011100000111101101000100100000010111001001"; --    +377325   +1181129
      WHEN  576 => Ti := "111111001011101111000110000011100110101010010111"; --    -214074    +944791
      WHEN  577 => Ti := "111100000101001011010010000000000101111011010101"; --   -1027374     +24277
      WHEN  578 => Ti := "000001010100101100111101111110111111100000010001"; --    +346941    -264175
      WHEN  579 => Ti := "000011001101111110101111000010011011100011011111"; --    +843695    +637151
      WHEN  580 => Ti := "000011110001100100001011000001010000100001101000"; --    +989451    +329832
      WHEN  581 => Ti := "111110111110110101110111111100011001110000001100"; --    -266889    -943092
      WHEN  582 => Ti := "000111100101000010010101000001011100000101011001"; --   +1986709    +377177
      WHEN  583 => Ti := "111110101010100011010010111001111100100100000010"; --    -349998   -1586942
      WHEN  584 => Ti := "000011001110001011100110000000111110010000101010"; --    +844518    +255018
      WHEN  585 => Ti := "000010011101000110010011000001011001110010010111"; --    +643475    +367767
      WHEN  586 => Ti := "000000011011010001111110000000010101111100111001"; --    +111742     +89913
      WHEN  587 => Ti := "000000100001000010010111000000111000100010101110"; --    +135319    +231598
      WHEN  588 => Ti := "111111111010010101101111000000110001100011110000"; --     -23185    +202992
      WHEN  589 => Ti := "111100010000000100100010111110000110110101011001"; --    -982750    -496295
      WHEN  590 => Ti := "000011101011101000010111000000000111111000001110"; --    +965143     +32270
      WHEN  591 => Ti := "000011000010000100010001000000000011101111000110"; --    +794897     +15302
      WHEN  592 => Ti := "000000011111011110100000000001110101011101011011"; --    +128928    +481115
      WHEN  593 => Ti := "000011101001100010000010000100010011111001001101"; --    +956546   +1130061
      WHEN  594 => Ti := "111011110110111010011011000000100110110101000110"; --   -1085797    +159046
      WHEN  595 => Ti := "111111110111000101011010111110000110010001011100"; --     -36518    -498596
      WHEN  596 => Ti := "000000100000010000110111000010000111011110010100"; --    +132151    +554900
      WHEN  597 => Ti := "000101010101100100010010000000101011000101111000"; --   +1399058    +176504
      WHEN  598 => Ti := "000000111110001011101101111111011011111010000001"; --    +254701    -147839
      WHEN  599 => Ti := "000001110000011110110100111110100000110000111100"; --    +460724    -390084
      WHEN  600 => Ti := "000100111110111110111101111110111100001100110001"; --   +1306557    -277711
      WHEN  601 => Ti := "111110001010110011011110111110010001111100100010"; --    -480034    -450782
      WHEN  602 => Ti := "111110011111111011111001000001100100010010001001"; --    -393479    +410761
      WHEN  603 => Ti := "000010101111100110110101000000000001011110011001"; --    +719285      +6041
      WHEN  604 => Ti := "000000100011101100010011111101001100000100011110"; --    +146195    -736994
      WHEN  605 => Ti := "000111010100111100000010111001111001110101010111"; --   +1920770   -1598121
      WHEN  606 => Ti := "000001110110010110111000000010011101000001110000"; --    +484792    +643184
      WHEN  607 => Ti := "111100011001101110111100000010001111100110110010"; --    -943172    +588210
      WHEN  608 => Ti := "111111101000110100011101111110000011000010000110"; --     -94947    -511866
      WHEN  609 => Ti := "111000111010101001001000111110001110001001011101"; --   -1856952    -466339
      WHEN  610 => Ti := "111100110001010100111100111111101111000000000000"; --    -846532     -69632
      WHEN  611 => Ti := "111101011001111001001010000011111001111011111100"; --    -680374   +1023740
      WHEN  612 => Ti := "111111111011110010100101000011001001110101101011"; --     -17243    +826731
      WHEN  613 => Ti := "000010110110111110111111000010001000100101011010"; --    +749503    +559450
      WHEN  614 => Ti := "000000101010111111010001000000001101111100010110"; --    +176081     +57110
      WHEN  615 => Ti := "000010010010111011100011000011000100000010010001"; --    +601827    +802961
      WHEN  616 => Ti := "111011111001000001000011000010000101111001101101"; --   -1077181    +548461
      WHEN  617 => Ti := "111101101100101000000111111101100001001001010111"; --    -603641    -650665
      WHEN  618 => Ti := "000000100001110001010110000100010110101111101100"; --    +138326   +1141740
      WHEN  619 => Ti := "000010101100010110100000111110101100011101011110"; --    +705952    -342178
      WHEN  620 => Ti := "000001001001110001001011111111100111000111011001"; --    +302155    -101927
      WHEN  621 => Ti := "000000000101001010100001000001000111010101100001"; --     +21153    +292193
      WHEN  622 => Ti := "000001110100010100100111000001100100110111100001"; --    +476455    +413153
      WHEN  623 => Ti := "111110111101100001110111000001010011001010111100"; --    -272265    +340668
      WHEN  624 => Ti := "111101000011001101110100111100110101100011111000"; --    -773260    -829192
      WHEN  625 => Ti := "111111011010011011000010111101100011011001010111"; --    -153918    -641449
      WHEN  626 => Ti := "000001100101010001101110111101110100110010100000"; --    +414830    -570208
      WHEN  627 => Ti := "111101001010011111000010111111100111001101010100"; --    -743486    -101548
      WHEN  628 => Ti := "111011011101011001110111000000111001100010000111"; --   -1190281    +235655
      WHEN  629 => Ti := "000000100100101100010100111111000001011110101000"; --    +150292    -256088
      WHEN  630 => Ti := "000100000110100000011011111101011110011001111000"; --   +1075227    -661896
      WHEN  631 => Ti := "000100001100111001001101000001110000100001011010"; --   +1101389    +460890
      WHEN  632 => Ti := "111111001110001111011111111011111110010000000101"; --    -203809   -1055739
      WHEN  633 => Ti := "000010100111011100000111000001111100100010100100"; --    +685831    +510116
      WHEN  634 => Ti := "111111110010110000000100000010011011010110100110"; --     -54268    +636326
      WHEN  635 => Ti := "111111011011001010110001000001010101001110101101"; --    -150863    +349101
      WHEN  636 => Ti := "111110101010000001101001000000010000110110011010"; --    -352151     +69018
      WHEN  637 => Ti := "111110010001111001001100111101111000011010110010"; --    -450996    -555342
      WHEN  638 => Ti := "111101101110101011000111000001000111111111010110"; --    -595257    +294870
      WHEN  639 => Ti := "000011000101100101011100111111000111111001000000"; --    +809308    -229824
      WHEN  640 => Ti := "111011110011111000101011111110010110110100100001"; --   -1098197    -430815
      WHEN  641 => Ti := "000100000111001100010101111110101011010000010110"; --   +1078037    -347114
      WHEN  642 => Ti := "000010001010000001110001111101110110001010110100"; --    +565361    -564556
      WHEN  643 => Ti := "000010100011001001111110111001010111001011001010"; --    +668286   -1740086
      WHEN  644 => Ti := "000011101110001111111100111111100000100000101010"; --    +975868    -128982
      WHEN  645 => Ti := "111100001101000101110011000010100010010011111110"; --    -994957    +664830
      WHEN  646 => Ti := "000000101111000111000011111101100101011101100100"; --    +192963    -632988
      WHEN  647 => Ti := "111010100010011011001111000001010100100110001110"; --   -1431857    +346510
      WHEN  648 => Ti := "111010110001010001111010111101011100110010111011"; --   -1371014    -668485
      WHEN  649 => Ti := "000011110100101000011001111101001011110110011001"; --   +1002009    -737895
      WHEN  650 => Ti := "111111001001010100101000000010001001111011001000"; --    -223960    +564936
      WHEN  651 => Ti := "111111010001111100000101111111101010001000001001"; --    -188667     -89591
      WHEN  652 => Ti := "111111000110110111001011000001111011011001111110"; --    -234037    +505470
      WHEN  653 => Ti := "111011111001110011010101111111010101111101100001"; --   -1073963    -172191
      WHEN  654 => Ti := "111110110000110101101110000000100100100010101100"; --    -324242    +149676
      WHEN  655 => Ti := "111101111011110100011001000000010101010110100110"; --    -541415     +87462
      WHEN  656 => Ti := "111111110000001111111011111110011001010111111110"; --     -64517    -420354
      WHEN  657 => Ti := "111111100101001110001000111111111110010000000111"; --    -109688      -7161
      WHEN  658 => Ti := "111110000001011110010000000001010001010101001100"; --    -518256    +333132
      WHEN  659 => Ti := "000011010010101010101001000010100101101000100110"; --    +862889    +678438
      WHEN  660 => Ti := "111100111000010011101001000100001011100001111100"; --    -817943   +1095804
      WHEN  661 => Ti := "000100001000111100100111000000101100010111000000"; --   +1085223    +181696
      WHEN  662 => Ti := "000010001011011011101010111111000010111011110110"; --    +571114    -250122
      WHEN  663 => Ti := "000001010000100010100100000001001101100101110110"; --    +329892    +317814
      WHEN  664 => Ti := "000000000011100000111000000000001010111100110011"; --     +14392     +44851
      WHEN  665 => Ti := "000000011110000000000001000010010101001100000011"; --    +122881    +611075
      WHEN  666 => Ti := "000010110001010011110100000001010101100110001011"; --    +726260    +350603
      WHEN  667 => Ti := "111111011111010100100000000010001001100011110100"; --    -133856    +563444
      WHEN  668 => Ti := "111110100110110011010011000011010100000111110110"; --    -365357    +868854
      WHEN  669 => Ti := "111111101100011011011100111111011110111000110011"; --     -80164    -135629
      WHEN  670 => Ti := "111111110001101000101010000110110010100001110011"; --     -58838   +1779827
      WHEN  671 => Ti := "111110101110100111101101111111111011010111000110"; --    -333331     -19002
      WHEN  672 => Ti := "111011111111101011101011000000010100111011001011"; --   -1049877     +85707
      WHEN  673 => Ti := "000101010100001101010001111101111111011110100101"; --   +1393489    -526427
      WHEN  674 => Ti := "111101111110011101001101000001000111000011011000"; --    -530611    +291032
      WHEN  675 => Ti := "000001000110110100111011111111111011110100010010"; --    +290107     -17134
      WHEN  676 => Ti := "111110001011001100000000111001001111010110011101"; --    -478464   -1772131
      WHEN  677 => Ti := "111111011111000001010000111010100011101100000110"; --    -135088   -1426682
      WHEN  678 => Ti := "111111011010000010111110000001101011000110011111"; --    -155458    +438687
      WHEN  679 => Ti := "111101001001001110100110111101100001101001000001"; --    -748634    -648639
      WHEN  680 => Ti := "111111100111110110011111111110010010001001110001"; --     -98913    -449935
      WHEN  681 => Ti := "000001000011101100001111111101110101000010100111"; --    +277263    -569177
      WHEN  682 => Ti := "000000100010000010001010111111111011010101101111"; --    +139402     -19089
      WHEN  683 => Ti := "000000111011111000001100111101010110101100011101"; --    +245260    -693475
      WHEN  684 => Ti := "111111110110010001101011111111101001010001111000"; --     -39829     -93064
      WHEN  685 => Ti := "000010100001010001100110111110001011000101011010"; --    +660582    -478886
      WHEN  686 => Ti := "000001100001101100011101111101100111111010111111"; --    +400157    -622913
      WHEN  687 => Ti := "111111001111111001001101111111110101000011110001"; --    -197043     -44815
      WHEN  688 => Ti := "111011000110110001000110111110010010110101101100"; --   -1283002    -447124
      WHEN  689 => Ti := "111110110101111110110001000001010011011101100010"; --    -303183    +341858
      WHEN  690 => Ti := "000001100011110001111101000001001011011110101111"; --    +408701    +309167
      WHEN  691 => Ti := "111111000001000111101111111101100000100001111111"; --    -257553    -653185
      WHEN  692 => Ti := "111101001111011001010011000001010001101010100001"; --    -723373    +334497
      WHEN  693 => Ti := "000010010001100010010101111111000001111101110000"; --    +596117    -254096
      WHEN  694 => Ti := "111111011001100110100100000000010010001100110111"; --    -157276     +74551
      WHEN  695 => Ti := "111110110010111101111111111111110110100011010000"; --    -315521     -38704
      WHEN  696 => Ti := "000110011000111011110101111111000100001010110001"; --   +1674997    -245071
      WHEN  697 => Ti := "111110100111010100000101000000101111101001100010"; --    -363259    +195170
      WHEN  698 => Ti := "000001011000000010011111000011001001010101101110"; --    +360607    +824686
      WHEN  699 => Ti := "000010110001110000011001111111001001111000110110"; --    +728089    -221642
      WHEN  700 => Ti := "111110000111101111100011000010011111110000011010"; --    -492573    +654362
      WHEN  701 => Ti := "000000110111011001110101000001100101010011000010"; --    +226933    +414914
      WHEN  702 => Ti := "111101101010001111101101000010110011101001010111"; --    -613395    +735831
      WHEN  703 => Ti := "000001010001001001101110111100000100011111110110"; --    +332398   -1030154
      WHEN  704 => Ti := "111111101110111100000100111101101010100001011101"; --     -69884    -612259
      WHEN  705 => Ti := "111111111010111100110010111101111001100011101001"; --     -20686    -550679
      WHEN  706 => Ti := "111100001010111001111111000001010100111010001010"; --   -1003905    +347786
      WHEN  707 => Ti := "000010101111111001001110111001111100101101101010"; --    +720462   -1586326
      WHEN  708 => Ti := "000011000111010110110011111101000100101000001100"; --    +816563    -767476
      WHEN  709 => Ti := "000010000111010011011110111111110110010000110101"; --    +554206     -39883
      WHEN  710 => Ti := "111111101111011110100010000100101110100011101011"; --     -67678   +1239275
      WHEN  711 => Ti := "000010110111001111001010000100100010001010000111"; --    +750538   +1188487
      WHEN  712 => Ti := "000100011011110101111011111111000010100011100111"; --   +1162619    -251673
      WHEN  713 => Ti := "000010010000100010111000000000101100001101111000"; --    +592056    +181112
      WHEN  714 => Ti := "000000010011101110001101111101101110101011010010"; --     +80781    -595246
      WHEN  715 => Ti := "000100011110111000100010111100110110001101100111"; --   +1175074    -826521
      WHEN  716 => Ti := "000011101101111100010110111110011110010111010111"; --    +974614    -399913
      WHEN  717 => Ti := "111111100001011010011101000011011100101010110001"; --    -125283    +903857
      WHEN  718 => Ti := "111110101010010000010011111111001100110111000010"; --    -351213    -209470
      WHEN  719 => Ti := "000001011001111110001111111111001011100100001100"; --    +368527    -214772
      WHEN  720 => Ti := "111110111100000011111010000000110010101111011000"; --    -278278    +207832
      WHEN  721 => Ti := "111111001101001100010001000001100111011101100100"; --    -208111    +423780
      WHEN  722 => Ti := "111110000110001110011101000101011110101100010000"; --    -498787   +1436432
      WHEN  723 => Ti := "111110111110011000111000111110101110010000011100"; --    -268744    -334820
      WHEN  724 => Ti := "111101011101000111110110111011110001111011101010"; --    -667146   -1106198
      WHEN  725 => Ti := "000000100001001001000001000000111000101100101000"; --    +135745    +232232
      WHEN  726 => Ti := "111100010100100000001000111101010100011010001100"; --    -964600    -702836
      WHEN  727 => Ti := "000000111101110101011111000000111010011010001100"; --    +253279    +239244
      WHEN  728 => Ti := "000010010000000000010110000011000001101010110110"; --    +589846    +793270
      WHEN  729 => Ti := "111111000110100111111100110110011111110111010100"; --    -235012   -2490924
      WHEN  730 => Ti := "000000001110010010000001111100110101100101010101"; --     +58497    -829099
      WHEN  731 => Ti := "111100010010110011010011000000001110010010100010"; --    -971565     +58530
      WHEN  732 => Ti := "111110011101001011000010111101010011101111100000"; --    -404798    -705568
      WHEN  733 => Ti := "111101010111010001111011000000001100110000110001"; --    -691077     +52273
      WHEN  734 => Ti := "111100010111111011010101000001011100100111100111"; --    -950571    +379367
      WHEN  735 => Ti := "000001100001010111110110111100111010011011111000"; --    +398838    -809224
      WHEN  736 => Ti := "000101101100110001001110000000001001110001010100"; --   +1494094     +40020
      WHEN  737 => Ti := "111100111001000010101101111100100010011010111110"; --    -814931    -907586
      WHEN  738 => Ti := "000001011100001011100110000000000110011111100001"; --    +377574     +26593
      WHEN  739 => Ti := "111011010010001000011101111101000011101111111000"; --   -1236451    -771080
      WHEN  740 => Ti := "000001100010011001110000111101111001000011001001"; --    +403056    -552759
      WHEN  741 => Ti := "111110111110100110010001000010111111011001001001"; --    -267887    +783945
      WHEN  742 => Ti := "000001001001100100011110000000001000000010111110"; --    +301342     +32958
      WHEN  743 => Ti := "111111111010110100000010111111010100101010110110"; --     -21246    -177482
      WHEN  744 => Ti := "000001010111000111110011111101101101001101101111"; --    +356851    -601233
      WHEN  745 => Ti := "000010001100010010000001111011000001101111011010"; --    +574593   -1303590
      WHEN  746 => Ti := "111100110010000100110000000000000110011100110000"; --    -843472     +26416
      WHEN  747 => Ti := "111101011011010100011011111100011010110100010001"; --    -674533    -938735
      WHEN  748 => Ti := "111111110001001111001000000000101001000000011010"; --     -60472    +167962
      WHEN  749 => Ti := "111111101101100011101001111011110101101101001111"; --     -75543   -1090737
      WHEN  750 => Ti := "000010000011000011001010000001001001001100101100"; --    +536778    +299820
      WHEN  751 => Ti := "000001001101100110010111000001011000100111001011"; --    +317847    +362955
      WHEN  752 => Ti := "000001111111110100101111000000100111100001110011"; --    +523567    +161907
      WHEN  753 => Ti := "111011101101001001101111000000101011010110101011"; --   -1125777    +177579
      WHEN  754 => Ti := "000010011111010010110111111111000000011100100101"; --    +652471    -260315
      WHEN  755 => Ti := "111110000100001000111101111111010000111111101111"; --    -507331    -192529
      WHEN  756 => Ti := "111101110110011010101101000000110001011010110000"; --    -563539    +202416
      WHEN  757 => Ti := "000000001001110001011001000011011001000000010111"; --     +40025    +888855
      WHEN  758 => Ti := "111111000110111100010111111100100011111001110000"; --    -233705    -901520
      WHEN  759 => Ti := "111111001101110001111111111101101110000100101000"; --    -205697    -597720
      WHEN  760 => Ti := "111010101110011010101111000000001110111000101100"; --   -1382737     +60972
      WHEN  761 => Ti := "111110001111101011110100000000010000100110000111"; --    -460044     +67975
      WHEN  762 => Ti := "000010110011010111100101000011010001100010000101"; --    +734693    +858245
      WHEN  763 => Ti := "000010100011000100001001111111111110110110100001"; --    +667913      -4703
      WHEN  764 => Ti := "111101101000110010010010111110101000011001101110"; --    -619374    -358802
      WHEN  765 => Ti := "111101100010011100000010111101110111000011110100"; --    -645374    -560908
      WHEN  766 => Ti := "000000110110100100101011000001101000001110001111"; --    +223531    +426895
      WHEN  767 => Ti := "000000001101111111111100000010000100110001111011"; --     +57340    +543867
      WHEN  768 => Ti := "000010110001001101101110000001110001001010001101"; --    +725870    +463501
      WHEN  769 => Ti := "000000101001001100111101000000011101101010101110"; --    +168765    +121518
      WHEN  770 => Ti := "000000011110010100010111111110110001001000110101"; --    +124183    -323019
      WHEN  771 => Ti := "000010000001010101011011111110001011010100001011"; --    +529755    -477941
      WHEN  772 => Ti := "000000000101000000011100000000001111010101001000"; --     +20508     +62792
      WHEN  773 => Ti := "000000010010100111000110111011001111011011010000"; --     +76230   -1247536
      WHEN  774 => Ti := "000100000001011111001100111100101000101001000101"; --   +1054668    -882107
      WHEN  775 => Ti := "111110001010011110000101000001010001010101001010"; --    -481403    +333130
      WHEN  776 => Ti := "000001000101110000111110111111010000000100010111"; --    +285758    -196329
      WHEN  777 => Ti := "000011000110101000100111111011111111101101101011"; --    +813607   -1049749
      WHEN  778 => Ti := "111111110011101000000010111111100111001010111001"; --     -50686    -101703
      WHEN  779 => Ti := "000011001100110011100101000010111010011111101001"; --    +838885    +763881
      WHEN  780 => Ti := "111101011000011111100000000000000111010111011010"; --    -686112     +30170
      WHEN  781 => Ti := "000100011001111010110101000010101000110100000111"; --   +1154741    +691463
      WHEN  782 => Ti := "111110100100001100100110000001100001101011110011"; --    -376026    +400115
      WHEN  783 => Ti := "111111101010011010001011000010101010100111101100"; --     -88437    +698860
      WHEN  784 => Ti := "000001000100001100100100000010101110101011000011"; --    +279332    +715459
      WHEN  785 => Ti := "111100000011000011000001111100011101111010101111"; --   -1036095    -926033
      WHEN  786 => Ti := "111111001000001110010111111111110011101111111011"; --    -228457     -50181
      WHEN  787 => Ti := "000001101011111011011011111101110000000001100110"; --    +442075    -589722
      WHEN  788 => Ti := "111010001100110100100101111110000100010011001110"; --   -1520347    -506674
      WHEN  789 => Ti := "111101110010111010011100000011100100001111100011"; --    -577892    +934883
      WHEN  790 => Ti := "000010000010011011111101111111000100100100011010"; --    +534269    -243430
      WHEN  791 => Ti := "111111000100111001010010111101100111101010110100"; --    -242094    -623948
      WHEN  792 => Ti := "111111001001000100101101000000011101001000001010"; --    -224979    +119306
      WHEN  793 => Ti := "000011001001111001101111000000110010110110011001"; --    +826991    +208281
      WHEN  794 => Ti := "111101111010010100000010000001110011110111101001"; --    -547582    +474601
      WHEN  795 => Ti := "111110101010100100100000000001100010101010110100"; --    -349920    +404148
      WHEN  796 => Ti := "000001001111110111111111000000111001010110001100"; --    +327167    +234892
      WHEN  797 => Ti := "111110101110100001111101111110101101011010010011"; --    -333699    -338285
      WHEN  798 => Ti := "111110000110110110010101000001100111000001100001"; --    -496235    +421985
      WHEN  799 => Ti := "111101101000000000000001111101110110011010100101"; --    -622591    -563547
      WHEN  800 => Ti := "111101111100101100011110111011110101110010001111"; --    -537826   -1090417
      WHEN  801 => Ti := "111011100101101011111111111111010011010010111100"; --   -1156353    -183108
      WHEN  802 => Ti := "111110101000000101110100111111001101100101010101"; --    -360076    -206507
      WHEN  803 => Ti := "111101010000101111011100111111110111111110010010"; --    -717860     -32878
      WHEN  804 => Ti := "000001110001111111110100111111101001111001010010"; --    +466932     -90542
      WHEN  805 => Ti := "111110011110001111111111000001011001110010011010"; --    -400385    +367770
      WHEN  806 => Ti := "000001000010111011101011000010011111101101011111"; --    +274155    +654175
      WHEN  807 => Ti := "000001110001110110111001000001010100100010001101"; --    +466361    +346253
      WHEN  808 => Ti := "000000100000011100110001000010100111010010001010"; --    +132913    +685194
      WHEN  809 => Ti := "000000111010111001011101111110110110100001101001"; --    +241245    -300951
      WHEN  810 => Ti := "111111111110011001011100000000011111110011010001"; --      -6564    +130257
      WHEN  811 => Ti := "111110010111100010100100000010100111110101001111"; --    -427868    +687439
      WHEN  812 => Ti := "111110100110010100000001111100111010100000000111"; --    -367359    -808953
      WHEN  813 => Ti := "111011011101110111000000111110010110100011000101"; --   -1188416    -431931
      WHEN  814 => Ti := "111101010100100101100000000100111001111000111110"; --    -702112   +1285694
      WHEN  815 => Ti := "111111100111101010101101000001000000100110010111"; --     -99667    +264599
      WHEN  816 => Ti := "111101000011010101010010111010000101110111111000"; --    -772782   -1548808
      WHEN  817 => Ti := "111110000111001001001100000100100011110001100110"; --    -495028   +1195110
      WHEN  818 => Ti := "111110000111011000111000000010011111011000100001"; --    -494024    +652833
      WHEN  819 => Ti := "111110111100010000101111000011011111111110101010"; --    -277457    +917418
      WHEN  820 => Ti := "111101100010111101101101000011000111011100110111"; --    -643219    +816951
      WHEN  821 => Ti := "000010100010110011101010000010110001100100010100"; --    +666858    +727316
      WHEN  822 => Ti := "000011001111000001000010000000100110011000111100"; --    +847938    +157244
      WHEN  823 => Ti := "000100010001000011101100000000011101111100100001"; --   +1118444    +122657
      WHEN  824 => Ti := "000101001100011010110110000001111101000010000010"; --   +1361590    +512130
      WHEN  825 => Ti := "111110101110001010111000111110010101110010111100"; --    -335176    -435012
      WHEN  826 => Ti := "111111110111101011101111111110111101101111001101"; --     -34065    -271411
      WHEN  827 => Ti := "111111000000000010110001111101000111010011100001"; --    -261967    -756511
      WHEN  828 => Ti := "000101000001111110111100000001001001011001001101"; --   +1318844    +300621
      WHEN  829 => Ti := "000010110001011110001011000001001011000001111101"; --    +726923    +307325
      WHEN  830 => Ti := "111111010111010101011110000010011100000001110000"; --    -166562    +639088
      WHEN  831 => Ti := "111111110101000110100100000001101100100100110011"; --     -44636    +444723
      WHEN  832 => Ti := "111111001001000111011001111110101001110111001000"; --    -224807    -352824
      WHEN  833 => Ti := "111111101001011110110101111111011110001001100010"; --     -92235    -138654
      WHEN  834 => Ti := "111111110010001010010100000011010100011010101101"; --     -56684    +870061
      WHEN  835 => Ti := "000000100010100011000010111110111101011110011001"; --    +141506    -272487
      WHEN  836 => Ti := "111110111000111101110100111110101010000001110000"; --    -290956    -352144
      WHEN  837 => Ti := "000011010110101011101010111110110001011010001000"; --    +879338    -321912
      WHEN  838 => Ti := "111100111000001001111010000001101110010000100001"; --    -818566    +451617
      WHEN  839 => Ti := "000001010111110111011001000010111101010100100000"; --    +359897    +775456
      WHEN  840 => Ti := "111110111001110110001100000101111101010110001101"; --    -287348   +1561997
      WHEN  841 => Ti := "000001101000101111011101000010101011001010111010"; --    +429021    +701114
      WHEN  842 => Ti := "000001101110111001011010000101100000111101101001"; --    +454234   +1445737
      WHEN  843 => Ti := "000010101111011101001101111110011111001010110101"; --    +718669    -396619
      WHEN  844 => Ti := "111110001110110111110111111110101101111000000000"; --    -463369    -336384
      WHEN  845 => Ti := "111111100100100111100011000000100001111110110011"; --    -112157    +139187
      WHEN  846 => Ti := "000001110010001000011110000101001100110111110011"; --    +467486   +1363443
      WHEN  847 => Ti := "111111100110000001100011111111001100000101110000"; --    -106397    -212624
      WHEN  848 => Ti := "111111000100111010111110000000011111100100011000"; --    -241986    +129304
      WHEN  849 => Ti := "000001001110000010110010000000111111010111101001"; --    +319666    +259561
      WHEN  850 => Ti := "000011100110010100000110000011010110110100011011"; --    +943366    +879899
      WHEN  851 => Ti := "000010011010100000000001111110100001000111001111"; --    +632833    -388657
      WHEN  852 => Ti := "111111110111110000001110111111101110001011000101"; --     -33778     -73019
      WHEN  853 => Ti := "111010011010011110111001000100101010011001111111"; --   -1464391   +1222271
      WHEN  854 => Ti := "111111100101010000001111000001010000011100001001"; --    -109553    +329481
      WHEN  855 => Ti := "000001010000011101000100000001011100011011111011"; --    +329540    +378619
      WHEN  856 => Ti := "000010001010001011100111111010111111001101110101"; --    +565991   -1313931
      WHEN  857 => Ti := "111010000111011010101011000000010110111100010101"; --   -1542485     +93973
      WHEN  858 => Ti := "111111111010001100110101000010011011011101110011"; --     -23755    +636787
      WHEN  859 => Ti := "111111101001110011101000000000001010111000111000"; --     -90904     +44600
      WHEN  860 => Ti := "000100111110111010101001111111011111001100000101"; --   +1306281    -134395
      WHEN  861 => Ti := "000101101010010110010110111011000101000110111111"; --   +1484182   -1289793
      WHEN  862 => Ti := "111111111110101010001111111101010011110111100110"; --      -5489    -705050
      WHEN  863 => Ti := "000011100111100001000110111101100101100001110101"; --    +948294    -632715
      WHEN  864 => Ti := "111111011111001000011010000010111001101011011110"; --    -134630    +760542
      WHEN  865 => Ti := "111101101111110000001010111101100010010101110000"; --    -590838    -645776
      WHEN  866 => Ti := "111110100101011100010111111011100010011001011101"; --    -370921   -1169827
      WHEN  867 => Ti := "111101111100101100011100111110011011000001011100"; --    -537828    -413604
      WHEN  868 => Ti := "000010000110000101001100111111101111100001001101"; --    +549196     -67507
      WHEN  869 => Ti := "000010101000101000011101000000100101000111111010"; --    +690717    +152058
      WHEN  870 => Ti := "000000010110111100111010000000100100110001101100"; --     +94010    +150636
      WHEN  871 => Ti := "000010010011100101100010111110101000000010001000"; --    +604514    -360312
      WHEN  872 => Ti := "000100011000101001110101000010010100000111101110"; --   +1149557    +606702
      WHEN  873 => Ti := "000010110000010101011000111100001001001100000100"; --    +722264   -1010940
      WHEN  874 => Ti := "000010010011100010111010111110010010111010100101"; --    +604346    -446811
      WHEN  875 => Ti := "111011110011000011110001000100010100000110001101"; --   -1101583   +1130893
      WHEN  876 => Ti := "000011101100000110011001000010000100000001111111"; --    +967065    +540799
      WHEN  877 => Ti := "111101011011110101000011111100001000001111100111"; --    -672445   -1014809
      WHEN  878 => Ti := "000011001101111101101110111101000001110100110000"; --    +843630    -778960
      WHEN  879 => Ti := "111110101010011000111011111100110101011101100011"; --    -350661    -829597
      WHEN  880 => Ti := "111111011101110110011011000000001100011001101011"; --    -139877     +50795
      WHEN  881 => Ti := "111101011000110111011010111111011110101001110001"; --    -684582    -136591
      WHEN  882 => Ti := "000000000110110010000011111110110100010111100100"; --     +27779    -309788
      WHEN  883 => Ti := "000001101111100111011111000011010101100100100111"; --    +457183    +874791
      WHEN  884 => Ti := "111010101101100010010000000000101001010100000101"; --   -1386352    +169221
      WHEN  885 => Ti := "111110100011000100101000000000000110000011100001"; --    -380632     +24801
      WHEN  886 => Ti := "111101100000001011011011000000101000010100111100"; --    -654629    +165180
      WHEN  887 => Ti := "111110110001101100110000000001011011100000011010"; --    -320720    +374810
      WHEN  888 => Ti := "000000011011110010010110000010101100100111011110"; --    +113814    +707038
      WHEN  889 => Ti := "111100011100101010100100111100111110111111000000"; --    -931164    -790592
      WHEN  890 => Ti := "111110101010101111111100000011110101000101010101"; --    -349188   +1003861
      WHEN  891 => Ti := "000000100111110110010111111101110111010000000011"; --    +163223    -560125
      WHEN  892 => Ti := "111101000100111011011110000101001000010101011001"; --    -766242   +1344857
      WHEN  893 => Ti := "111110101000000101001110111110011110010111010010"; --    -360114    -399918
      WHEN  894 => Ti := "111111000101110111111001000001101000111001111100"; --    -238087    +429692
      WHEN  895 => Ti := "000001001011010110110010000000100000011011001111"; --    +308658    +132815
      WHEN  896 => Ti := "000011001000101010001100111110010011101001000101"; --    +821900    -443835
      WHEN  897 => Ti := "000000001100110100110001111110010000001110011000"; --     +52529    -457832
      WHEN  898 => Ti := "111110000001101000001100000000111111010011101110"; --    -517620    +259310
      WHEN  899 => Ti := "000011110000111001000100000001111101100001101100"; --    +986692    +514156
      WHEN  900 => Ti := "000001101011111001111010000011000111111001010001"; --    +441978    +818769
      WHEN  901 => Ti := "000000000011011000111010111111100111011000001010"; --     +13882    -100854
      WHEN  902 => Ti := "111110110001010010111111111100111101111010110111"; --    -322369    -794953
      WHEN  903 => Ti := "000000110111000100011000000001011010100011101010"; --    +225560    +370922
      WHEN  904 => Ti := "000000000001110110100100000001111100001001010101"; --      +7588    +508501
      WHEN  905 => Ti := "000010011011100100110011111101110001111010101000"; --    +637235    -581976
      WHEN  906 => Ti := "000000101010000100110111111110000100010100101001"; --    +172343    -506583
      WHEN  907 => Ti := "000001001010101011010101000000000110001110000000"; --    +305877     +25472
      WHEN  908 => Ti := "000001101001010001000101000001011100101010101000"; --    +431173    +379560
      WHEN  909 => Ti := "000010011111111100110111000011101011110111011010"; --    +655159    +966106
      WHEN  910 => Ti := "000101010001100011011001111111100111111100000011"; --   +1382617     -98557
      WHEN  911 => Ti := "111100101110010010101100000001001011011000111000"; --    -858964    +308792
      WHEN  912 => Ti := "000001100101011100011000111111000001010100101111"; --    +415512    -256721
      WHEN  913 => Ti := "000100000001010101001001000010000000110010110110"; --   +1054025    +527542
      WHEN  914 => Ti := "000001101001011000011001000100010101000111110010"; --    +431641   +1135090
      WHEN  915 => Ti := "000001010000000000101011111011110111111010101001"; --    +327723   -1081687
      WHEN  916 => Ti := "111111001010111001000010000011000000111010101100"; --    -217534    +790188
      WHEN  917 => Ti := "000001011000010110010111000000101110000010000100"; --    +361879    +188548
      WHEN  918 => Ti := "111111000010111000101010111110111000000101011111"; --    -250326    -294561
      WHEN  919 => Ti := "111100000011100000110000111111101100010110110111"; --   -1034192     -80457
      WHEN  920 => Ti := "000000011001110110001000000001001000011110011000"; --    +105864    +296856
      WHEN  921 => Ti := "000000111001111100111100111110000000111011101111"; --    +237372    -520465
      WHEN  922 => Ti := "111111100110111010100010000000001110111101101111"; --    -102750     +61295
      WHEN  923 => Ti := "000001110101010000110001000001010011011110000110"; --    +480305    +341894
      WHEN  924 => Ti := "111110101000101000010001000100000101000000111100"; --    -357871   +1069116
      WHEN  925 => Ti := "000000001000110000010101111111011000001010011110"; --     +35861    -163170
      WHEN  926 => Ti := "000000011101101000101100111111000101010101001001"; --    +121388    -240311
      WHEN  927 => Ti := "000000010111100110011100111010100010011101101011"; --     +96668   -1431701
      WHEN  928 => Ti := "000001100100110010011010111111000011000111111101"; --    +412826    -249347
      WHEN  929 => Ti := "111111000011100000101010111111011111101001100111"; --    -247766    -132505
      WHEN  930 => Ti := "111101010010110100101100000000111000111101110110"; --    -709332    +233334
      WHEN  931 => Ti := "000101010001001111000000111101111001011000001011"; --   +1381312    -551413
      WHEN  932 => Ti := "000001011011001001111001111101011100100000101100"; --    +373369    -669652
      WHEN  933 => Ti := "000011001111100101000001000001000110000101111001"; --    +850241    +287097
      WHEN  934 => Ti := "111110000110011111101011111110101001100110101110"; --    -497685    -353874
      WHEN  935 => Ti := "000000111100110101001111111101110000011001100001"; --    +249167    -588191
      WHEN  936 => Ti := "111111101101111000101010000000011101010011110001"; --     -74198    +120049
      WHEN  937 => Ti := "111011111011001001011001111001011010011001100111"; --   -1068455   -1726873
      WHEN  938 => Ti := "000000000100110100011100000100100001110101001100"; --     +19740   +1187148
      WHEN  939 => Ti := "111010100000001100100011111111110100100110101111"; --   -1440989     -46673
      WHEN  940 => Ti := "000011110110111001000000000000000010000101111000"; --   +1011264      +8568
      WHEN  941 => Ti := "111110100111101101101001111011000001101110100101"; --    -361623   -1303643
      WHEN  942 => Ti := "111100111111100101111111000001010001001001001110"; --    -788097    +332366
      WHEN  943 => Ti := "111111000111000011111100000000010011111000100001"; --    -233220     +81441
      WHEN  944 => Ti := "111111111111110000100110111100100111111010110100"; --       -986    -885068
      WHEN  945 => Ti := "000011001101111101011110000001010100110100111000"; --    +843614    +347448
      WHEN  946 => Ti := "111111000010101010000111111111011011110110110010"; --    -251257    -148046
      WHEN  947 => Ti := "111100101000011011100000111101100000110011010100"; --    -882976    -652076
      WHEN  948 => Ti := "111100000001111011001101111101101000011001001001"; --   -1040691    -620983
      WHEN  949 => Ti := "111100000111000101011101000000011001011111101111"; --   -1019555    +104431
      WHEN  950 => Ti := "000001000010001001110110111101100101101011000000"; --    +270966    -632128
      WHEN  951 => Ti := "000011010110000011111111111101101011100010111011"; --    +876799    -608069
      WHEN  952 => Ti := "111100101101111111011101111110110110110100110111"; --    -860195    -299721
      WHEN  953 => Ti := "111111011101111100111101111101100011111101110101"; --    -139459    -639115
      WHEN  954 => Ti := "000001000100110001101100000010001010010100111100"; --    +281708    +566588
      WHEN  955 => Ti := "000010011101011111101000000010010111000000101101"; --    +645096    +618541
      WHEN  956 => Ti := "111110000001000000000001111110010101000110010011"; --    -520191    -437869
      WHEN  957 => Ti := "111111010111111100010101000000010110110101100111"; --    -164075     +93543
      WHEN  958 => Ti := "111000010011010100101111110111111011010000001011"; --   -2018001   -2116597
      WHEN  959 => Ti := "000001011011100011110101111101100011001100101111"; --    +375029    -642257
      WHEN  960 => Ti := "111110000110100001101001111111110001111011011101"; --    -497559     -57635
      WHEN  961 => Ti := "000010101111101110011110111111100111011000110011"; --    +719774    -100813
      WHEN  962 => Ti := "000000000101110001001101000010000101011101100111"; --     +23629    +546663
      WHEN  963 => Ti := "000001000011111101010100111101011111011001000111"; --    +278356    -657849
      WHEN  964 => Ti := "111101110001101001111110000001000101100000110010"; --    -583042    +284722
      WHEN  965 => Ti := "111001101101011100111100000010001010011001000101"; --   -1648836    +566853
      WHEN  966 => Ti := "111111100111101111111111000010011001110101101011"; --     -99329    +630123
      WHEN  967 => Ti := "000001000101010000100111111110100110001001000101"; --    +283687    -368059
      WHEN  968 => Ti := "000000010001101000011000111110000010100011101101"; --     +72216    -513811
      WHEN  969 => Ti := "000001000011110101110001111011010100110010100000"; --    +277873   -1225568
      WHEN  970 => Ti := "111110000010001011101011000001001011010111110011"; --    -515349    +308723
      WHEN  971 => Ti := "000000100011101101001111000001000111101011001100"; --    +146255    +293580
      WHEN  972 => Ti := "111011111110010100000010111110001110000100010010"; --   -1055486    -466670
      WHEN  973 => Ti := "111110001000010100010010111111110110000010001100"; --    -490222     -40820
      WHEN  974 => Ti := "000100111100100111000010000010010111110001001100"; --   +1296834    +621644
      WHEN  975 => Ti := "111111101001000110100101000000010101100001111110"; --     -93787     +88190
      WHEN  976 => Ti := "000010011011011011111101000100111100001100101100"; --    +636669   +1295148
      WHEN  977 => Ti := "111110110110001111010001000001100010100110001101"; --    -302127    +403853
      WHEN  978 => Ti := "000010111101110100001110111110011011111011100111"; --    +777486    -409881
      WHEN  979 => Ti := "000001111000000000111111000011101010010011111001"; --    +491583    +959737
      WHEN  980 => Ti := "000001001010111110000110000010101001000101111111"; --    +307078    +692607
      WHEN  981 => Ti := "111111001100000010111000000000011101011100101101"; --    -212808    +120621
      WHEN  982 => Ti := "111101010101101011010100111110110110101010111010"; --    -697644    -300358
      WHEN  983 => Ti := "000010010000000101001101000000001101101110010011"; --    +590157     +56211
      WHEN  984 => Ti := "111111110100001000110111000111000100101001111110"; --     -48585   +1854078
      WHEN  985 => Ti := "111110100111111001000111111011111010111001000010"; --    -360889   -1069502
      WHEN  986 => Ti := "000000111000001001000010111110101110001000011101"; --    +229954    -335331
      WHEN  987 => Ti := "000000111011101010111111000100010110111111000110"; --    +244415   +1142726
      WHEN  988 => Ti := "111100111001001101110111000001111010100000000010"; --    -814217    +501762
      WHEN  989 => Ti := "111110011001001111101011111111111101001001100001"; --    -420885     -11679
      WHEN  990 => Ti := "000011011100100101010001000001100010110111001110"; --    +903505    +404942
      WHEN  991 => Ti := "000000111011100001000111000000111111110110110110"; --    +243783    +261558
      WHEN  992 => Ti := "111111000111000011001111000001000110000100000100"; --    -233265    +286980
      WHEN  993 => Ti := "000000000010011100011101111111000001101101001100"; --     +10013    -255156
      WHEN  994 => Ti := "111110010101110011110111000101000100110000011111"; --    -434953   +1330207
      WHEN  995 => Ti := "000100101110101100100011000010100001001010100101"; --   +1239843    +660133
      WHEN  996 => Ti := "111110000001100101110010111101100100110111001100"; --    -517774    -635444
      WHEN  997 => Ti := "111101000111111000100110000111101101111101111010"; --    -754138   +2023290
      WHEN  998 => Ti := "111110111100101100100110000001010001100001110001"; --    -275674    +333937
      WHEN  999 => Ti := "111110011000111110111100111101110110001011111001"; --    -421956    -564487
      WHEN 1000 => Ti := "000001010000110100110101111110100100110011100110"; --    +331061    -373530
      WHEN 1001 => Ti := "000000010001110011111101000001011111111011000111"; --     +72957    +392903
      WHEN 1002 => Ti := "000110010001100110011010111110101011010001101011"; --   +1644954    -347029
      WHEN 1003 => Ti := "000010000010101001011010111111011010001101001100"; --    +535130    -154804
      WHEN 1004 => Ti := "111100110100001110110111111110010101001101101101"; --    -834633    -437395
      WHEN 1005 => Ti := "111110000110010100011011000010111100001100101100"; --    -498405    +770860
      WHEN 1006 => Ti := "000010100001011111111011000000101101110101101100"; --    +661499    +187756
      WHEN 1007 => Ti := "000000000110110000111001000100011101000111000000"; --     +27705   +1167808
      WHEN 1008 => Ti := "111011011111011001111000000100000101001110010100"; --   -1182088   +1069972
      WHEN 1009 => Ti := "111110110100111110110010111110111100100000100101"; --    -307278    -276443
      WHEN 1010 => Ti := "111111000010110101101111111110101010010010001010"; --    -250513    -351094
      WHEN 1011 => Ti := "000001000101000111001011111101111001111001100010"; --    +283083    -549278
      WHEN 1012 => Ti := "111111001011100011000101111101110010100000101110"; --    -214843    -579538
      WHEN 1013 => Ti := "000110000110001001110011000000001011010111001010"; --   +1598067     +46538
      WHEN 1014 => Ti := "000100010010001011001000000010001010111010010101"; --   +1123016    +568981
      WHEN 1015 => Ti := "000010100100010110010110000000010100111001100000"; --    +673174     +85600
      WHEN 1016 => Ti := "111001110010100110101011000010110001110010110000"; --   -1627733    +728240
      WHEN 1017 => Ti := "000001100000001100111101111110111000000001100110"; --    +394045    -294810
      WHEN 1018 => Ti := "000000001110111100010000111110101101011010000111"; --     +61200    -338297
      WHEN 1019 => Ti := "111110001110000011100001000001011011000000110000"; --    -466719    +372784
      WHEN 1020 => Ti := "000011011110100100001001111101101010111000100111"; --    +911625    -610777
      WHEN 1021 => Ti := "000010001000110111000100000001110111100110101111"; --    +560580    +489903
      WHEN 1022 => Ti := "111110010001111001000100000010001000101000110000"; --    -451004    +559664
      WHEN 1023 => Ti := "000001110010011011000001000000010000010100001001"; --    +468673     +66825
      WHEN 1024 => Ti := "000100111100111100100010000111001111001011011001"; --   +1298210   +1897177
      WHEN 1025 => Ti := "111111110101101111100001111110000111010110110101"; --     -42015    -494155
      WHEN 1026 => Ti := "000010111110001011011010000010110011011001010011"; --    +778970    +734803
      WHEN 1027 => Ti := "111100100011110101010001000001000010001111100100"; --    -901807    +271332
      WHEN 1028 => Ti := "000000111111110001110001111100111101001111001110"; --    +261233    -797746
      WHEN 1029 => Ti := "111101010110111011101000000100111001000101001101"; --    -692504   +1282381
      WHEN 1030 => Ti := "111100110100101111100110000001011100000101111111"; --    -832538    +377215
      WHEN 1031 => Ti := "000000101111000010101111111101010011011110001100"; --    +192687    -706676
      WHEN 1032 => Ti := "000011101000010110101010000010011001000010101111"; --    +951722    +626863
      WHEN 1033 => Ti := "000100011101100101100000000001010010001111000101"; --   +1169760    +336837
      WHEN 1034 => Ti := "111111000100101100100111111110111111000010010000"; --    -242905    -266096
      WHEN 1035 => Ti := "111100101011001111010101111100000100011010100101"; --    -871467   -1030491
      WHEN 1036 => Ti := "111111000000010001000001000100011110001001011010"; --    -261055   +1172058
      WHEN 1037 => Ti := "000000001111010000001101000011111001001100100011"; --     +62477   +1020707
      WHEN 1038 => Ti := "000001011100111110111100000001011101001100010010"; --    +380860    +381714
      WHEN 1039 => Ti := "111011010110101101110100000001100000001010111111"; --   -1217676    +393919
      WHEN 1040 => Ti := "111110011010011100100011111111000100111101000000"; --    -415965    -241856
      WHEN 1041 => Ti := "000001100001110010011101111110000110011101101010"; --    +400541    -497814
      WHEN 1042 => Ti := "000011011001100100001111000000111000001010101000"; --    +891151    +230056
      WHEN 1043 => Ti := "111111001100110001100111111111011111001110101110"; --    -209817    -134226
      WHEN 1044 => Ti := "111111100001010100111000000010010100011011000001"; --    -125640    +607937
      WHEN 1045 => Ti := "111110001000101100001110000000010010101111100011"; --    -488690     +76771
      WHEN 1046 => Ti := "000001000110000110000001000011000011010010000110"; --    +287105    +799878
      WHEN 1047 => Ti := "000000001100011010110100111001011001010011010111"; --     +50868   -1731369
      WHEN 1048 => Ti := "000001110110110010011110000000001110010110010001"; --    +486558     +58769
      WHEN 1049 => Ti := "000010010001010000011111000001110111100011000011"; --    +594975    +489667
      WHEN 1050 => Ti := "111110101101100100010101000001101101100010111001"; --    -337643    +448697
      WHEN 1051 => Ti := "111110001100101010111111000101000101111100100110"; --    -472385   +1335078
      WHEN 1052 => Ti := "000011001110011000100010000000110011101000110000"; --    +845346    +211504
      WHEN 1053 => Ti := "000000011011110111001010111101100010110011010100"; --    +114122    -643884
      WHEN 1054 => Ti := "111110111101000011101111000001010111100100011111"; --    -274193    +358687
      WHEN 1055 => Ti := "000011011001110001110010000001001010000101000010"; --    +892018    +303426
      WHEN 1056 => Ti := "111110010101100101000110000001001000110000010110"; --    -435898    +298006
      WHEN 1057 => Ti := "111100010010010110011110111010110001000110110101"; --    -973410   -1371723
      WHEN 1058 => Ti := "111111000101110001100111111110000100110111111001"; --    -238489    -504327
      WHEN 1059 => Ti := "000000010000001010011000000000001111101100000010"; --     +66200     +64258
      WHEN 1060 => Ti := "000001111100100111100101000011110100010001011100"; --    +510437   +1000540
      WHEN 1061 => Ti := "111101001100110010111110000100000111110001001110"; --    -734018   +1080398
      WHEN 1062 => Ti := "000100010001101011100010000001000000010011010101"; --   +1120994    +263381
      WHEN 1063 => Ti := "111101011101011011010101111110010010001110011010"; --    -665899    -449638
      WHEN 1064 => Ti := "111110011010010110001011000101010111001001111001"; --    -416373   +1405561
      WHEN 1065 => Ti := "111101101111011001101100000011010111101001110010"; --    -592276    +883314
      WHEN 1066 => Ti := "111100001000011100000001000000110001000110111000"; --   -1014015    +201144
      WHEN 1067 => Ti := "111110011110000011101011000011000110111001010101"; --    -401173    +814677
      WHEN 1068 => Ti := "111101010110001001111011000001000111100010101011"; --    -695685    +293035
      WHEN 1069 => Ti := "111101100011101110000111000100010011000101011001"; --    -640121   +1126745
      WHEN 1070 => Ti := "000001101010000110111100000100110110011011101010"; --    +434620   +1271530
      WHEN 1071 => Ti := "000010001110011101110110111111001011000010010110"; --    +583542    -216938
      WHEN 1072 => Ti := "111111001010000010100111000000001000111001111101"; --    -221017     +36477
      WHEN 1073 => Ti := "111111111111110111100111111101000010100111011111"; --       -537    -775713
      WHEN 1074 => Ti := "000100010110000101000001111111010011110000001010"; --   +1139009    -181238
      WHEN 1075 => Ti := "111110001110010011111101111100100110111001111000"; --    -465667    -889224
      WHEN 1076 => Ti := "111111110100011110000010111010011111000110111101"; --     -47230   -1445443
      WHEN 1077 => Ti := "111010101001111100110000000010100010010111101011"; --   -1401040    +665067
      WHEN 1078 => Ti := "000010010101001101110010111101010111001011010111"; --    +611186    -691497
      WHEN 1079 => Ti := "111110000001111110011010111000100001010101000000"; --    -516198   -1960640
      WHEN 1080 => Ti := "111010110011100000101101111111001101010101110111"; --   -1361875    -207497
      WHEN 1081 => Ti := "000101000111010110110011111100010111110100100101"; --   +1340851    -951003
      WHEN 1082 => Ti := "000000111111010000011101111111000001110001000001"; --    +259101    -254911
      WHEN 1083 => Ti := "000000000101010100010111111110001011000000000011"; --     +21783    -479229
      WHEN 1084 => Ti := "000000010011001111010110000000000110011101011000"; --     +78806     +26456
      WHEN 1085 => Ti := "000010100111010001001111000001100010011010111001"; --    +685135    +403129
      WHEN 1086 => Ti := "111110110001011111101001000100101101101000110101"; --    -321559   +1235509
      WHEN 1087 => Ti := "000000011010011010011000111110001000001101010110"; --    +108184    -490666
      WHEN 1088 => Ti := "111111010010111111110111000000011101000010110000"; --    -184329    +118960
      WHEN 1089 => Ti := "111111100110111111011111000001011111011101011100"; --    -102433    +391004
      WHEN 1090 => Ti := "000100100100101111100010000001100001111101010111"; --   +1199074    +401239
      WHEN 1091 => Ti := "000001111100000100011000111110111100001101001100"; --    +508184    -277684
      WHEN 1092 => Ti := "000001010101011100100110111110101101010110011000"; --    +349990    -338536
      WHEN 1093 => Ti := "000100110011001000000111000010111101100110001111"; --   +1257991    +776591
      WHEN 1094 => Ti := "111111110000111000101111000000111000010001010100"; --     -61905    +230484
      WHEN 1095 => Ti := "000010001110000011111001000010000100011011011011"; --    +581881    +542427
      WHEN 1096 => Ti := "111011001011100000001111111011111010001110101101"; --   -1263601   -1072211
      WHEN 1097 => Ti := "000001000101111111111100000001001101101101010101"; --    +286716    +318293
      WHEN 1098 => Ti := "111110110010001010010010111111110011110101000110"; --    -318830     -49850
      WHEN 1099 => Ti := "000000111100111011010011000000000010100011100110"; --    +249555     +10470
      WHEN 1100 => Ti := "000010100110001110110111111100000110010011010000"; --    +680887   -1022768
      WHEN 1101 => Ti := "111111001110111111011001000001010111011100101000"; --    -200743    +358184
      WHEN 1102 => Ti := "111101000000101000110001000001100111101001100110"; --    -783823    +424550
      WHEN 1103 => Ti := "000000001011011111111010000010101101111001011101"; --     +47098    +712285
      WHEN 1104 => Ti := "000000000110010001100100111110111111001110100001"; --     +25700    -265311
      WHEN 1105 => Ti := "111110000110011110011011111111101100010010100101"; --    -497765     -80731
      WHEN 1106 => Ti := "111100011000000101101100000010010010101001100110"; --    -949908    +600678
      WHEN 1107 => Ti := "000000101101011000010000000000001010011000010001"; --    +185872     +42513
      WHEN 1108 => Ti := "111110100111101110101101111010011110000101111010"; --    -361555   -1449606
      WHEN 1109 => Ti := "111101000101110110001111111101110110101111001000"; --    -762481    -562232
      WHEN 1110 => Ti := "111110010011110100110110111111001001010110100111"; --    -443082    -223833
      WHEN 1111 => Ti := "111111111111010111011111000011000010101101111000"; --      -2593    +797560
      WHEN 1112 => Ti := "000000000111011111000000000000101111100000011001"; --     +30656    +194585
      WHEN 1113 => Ti := "111101001010001010111011000010000110010111110111"; --    -744773    +550391
      WHEN 1114 => Ti := "000000001100011011111000111111101111000010111111"; --     +50936     -69441
      WHEN 1115 => Ti := "000000110010100000001101000001110011011110110001"; --    +206861    +473009
      WHEN 1116 => Ti := "000010011001111100011100000011011010111010101111"; --    +630556    +896687
      WHEN 1117 => Ti := "111101111010001001011100111111100000101110101000"; --    -548260    -128088
      WHEN 1118 => Ti := "000011110011101110000111111101011001111100000010"; --    +998279    -680190
      WHEN 1119 => Ti := "111101001001110000011001000010110000001010010000"; --    -746471    +721552
      WHEN 1120 => Ti := "000001100100010110110001111111110110100010110100"; --    +411057     -38732
      WHEN 1121 => Ti := "111010100010101100001111000000111011100101110010"; --   -1430769    +244082
      WHEN 1122 => Ti := "000010100101010101001010000000000010001101101010"; --    +677194      +9066
      WHEN 1123 => Ti := "111111110000110001001011111100001101100010001101"; --     -62389    -993139
      WHEN 1124 => Ti := "111100000011101110111111111100110100100100010100"; --   -1033281    -833260
      WHEN 1125 => Ti := "111110010000101110001010000000011100001100001100"; --    -455798    +115468
      WHEN 1126 => Ti := "111110010000011001010100000100101011110101010011"; --    -457132   +1228115
      WHEN 1127 => Ti := "000001010100101001100111111101010110101000101101"; --    +346727    -693715
      WHEN 1128 => Ti := "000010110000011101111110000100001110001011110101"; --    +722814   +1106677
      WHEN 1129 => Ti := "000101000000101110110100000000110001011100110011"; --   +1313716    +202547
      WHEN 1130 => Ti := "111111110001110100111110111110111000111100110011"; --     -58050    -291021
      WHEN 1131 => Ti := "111111010011111111110100111011111000101001001000"; --    -180236   -1078712
      WHEN 1132 => Ti := "000001001101001110110000111101011010101001111010"; --    +316336    -677254
      WHEN 1133 => Ti := "111100010010001001101011111110100110000100010001"; --    -974229    -368367
      WHEN 1134 => Ti := "000011111101001101111011000101000101111011110111"; --   +1037179   +1335031
      WHEN 1135 => Ti := "111111110100101101010000000001000001110101100110"; --     -46256    +269670
      WHEN 1136 => Ti := "111011101101001111111010111100000010011110111101"; --   -1125382   -1038403
      WHEN 1137 => Ti := "111100011011010010101100000010010111111101100000"; --    -936788    +622432
      WHEN 1138 => Ti := "111110101001000001001101000011111100000100100001"; --    -356275   +1032481
      WHEN 1139 => Ti := "111110110010001011100100000000010000101010000011"; --    -318748     +68227
      WHEN 1140 => Ti := "111111100111111111100010000011101100100000011111"; --     -98334    +968735
      WHEN 1141 => Ti := "111110111001000101100111000010000100111110000010"; --    -290457    +544642
      WHEN 1142 => Ti := "111111101101100101000010111111101010101000110110"; --     -75454     -87498
      WHEN 1143 => Ti := "111111011011010010000111111011110011000001001011"; --    -150393   -1101749
      WHEN 1144 => Ti := "111101011111011001011001111111011010010011010011"; --    -657831    -154413
      WHEN 1145 => Ti := "000001101100001101101101111111011000111110101010"; --    +443245    -159830
      WHEN 1146 => Ti := "000100001111010100011000000010000110001010011100"; --   +1111320    +549532
      WHEN 1147 => Ti := "000001001101110101010110111101010001100111101110"; --    +318806    -714258
      WHEN 1148 => Ti := "111110001011101001101111111110000001110011010001"; --    -476561    -516911
      WHEN 1149 => Ti := "111111000010100110110100111110000100011110000100"; --    -251468    -505980
      WHEN 1150 => Ti := "000100100101111101111011111011011010011101000100"; --   +1204091   -1202364
      WHEN 1151 => Ti := "000000011110101101010001111111110110010011001101"; --    +125777     -39731
      WHEN 1152 => Ti := "111111000111100000000010111111000110111000000100"; --    -231422    -233980
      WHEN 1153 => Ti := "000001001110010011110110111001111101111011101110"; --    +320758   -1581330
      WHEN 1154 => Ti := "000001101110000010110011000010110111101011001011"; --    +450739    +752331
      WHEN 1155 => Ti := "000010000101100000101000000010011100001010000000"; --    +546856    +639616
      WHEN 1156 => Ti := "111010100000101010100100111110001010101100101011"; --   -1439068    -480469
      WHEN 1157 => Ti := "111101110111110111001101111111100101111100010110"; --    -557619    -106730
      WHEN 1158 => Ti := "111111011010101001000010111110110110101111000000"; --    -153022    -300096
      WHEN 1159 => Ti := "111111101001100010110011000001111111101000101010"; --     -91981    +522794
      WHEN 1160 => Ti := "111110111110111011111111111101110001010110011100"; --    -266497    -584292
      WHEN 1161 => Ti := "000001001111101001001001000010110000110001011100"; --    +326217    +724060
      WHEN 1162 => Ti := "000011001111111001010000000010011011110011001111"; --    +851536    +638159
      WHEN 1163 => Ti := "111100101001110011101000111101101111110000101100"; --    -877336    -590804
      WHEN 1164 => Ti := "000001111000111001011101111110111101011100111000"; --    +495197    -272584
      WHEN 1165 => Ti := "111110011011110110110101000011000000111001101110"; --    -410187    +790126
      WHEN 1166 => Ti := "111100100000011110011111000010001101011011100001"; --    -915553    +579297
      WHEN 1167 => Ti := "111111111111000100000001111011100011011001110111"; --      -3839   -1165705
      WHEN 1168 => Ti := "111100111001001100011011111111001010001101001111"; --    -814309    -220337
      WHEN 1169 => Ti := "111111101101010010110010000001001101100110000011"; --     -76622    +317827
      WHEN 1170 => Ti := "000010100000010010101000111100101110001001100101"; --    +656552    -859547
      WHEN 1171 => Ti := "000010011010010000001001111111010110101110000101"; --    +631817    -169083
      WHEN 1172 => Ti := "111111000111010001001101000011110100000101100110"; --    -232371    +999782
      WHEN 1173 => Ti := "111111000010011000101011111110100011011101111010"; --    -252373    -379014
      WHEN 1174 => Ti := "111110101010010011100000000000100011110000011011"; --    -351008    +146459
      WHEN 1175 => Ti := "000000101100011111000010111101100000011111111111"; --    +182210    -653313
      WHEN 1176 => Ti := "000010001100011100111100000000101110110001010000"; --    +575292    +191568
      WHEN 1177 => Ti := "111101111100110001111011111110010001110001111110"; --    -537477    -451458
      WHEN 1178 => Ti := "000001101000101101111000111111101111011100010101"; --    +428920     -67819
      WHEN 1179 => Ti := "111101101011010100100101111110110110101111111010"; --    -608987    -300038
      WHEN 1180 => Ti := "111110110001100010111110000010110100111001110100"; --    -321346    +740980
      WHEN 1181 => Ti := "000101000101011001110000000010001010110101011101"; --   +1332848    +568669
      WHEN 1182 => Ti := "111110111110001011101010111111110101100101000111"; --    -269590     -42681
      WHEN 1183 => Ti := "000100001111111110010010000000000110101100011111"; --   +1114002     +27423
      WHEN 1184 => Ti := "111111100101101101010010111110010100000000001000"; --    -107694    -442360
      WHEN 1185 => Ti := "000010010010111100000000000001110110111110010100"; --    +601856    +487316
      WHEN 1186 => Ti := "111010110110011110011110000001101010100011000000"; --   -1349730    +436416
      WHEN 1187 => Ti := "000001110110101110000111111001100111001011010000"; --    +486279   -1674544
      WHEN 1188 => Ti := "111101001001110111010101000001100110111011111110"; --    -746027    +421630
      WHEN 1189 => Ti := "111101001011110010110001000000010000000101111010"; --    -738127     +65914
      WHEN 1190 => Ti := "111010100111001010101011000011010011110100010001"; --   -1412437    +867601
      WHEN 1191 => Ti := "000011011001101010110001111101100110010111010011"; --    +891569    -629293
      WHEN 1192 => Ti := "000000001000111100000100111110000001010001111110"; --     +36612    -519042
      WHEN 1193 => Ti := "000000011110100011110111111100011001011011111011"; --    +125175    -944389
      WHEN 1194 => Ti := "111100111111001111010110111101010101011001000000"; --    -789546    -698816
      WHEN 1195 => Ti := "111101001010011000011110111110101010001101000100"; --    -743906    -351420
      WHEN 1196 => Ti := "000000110111011000111011111110111111110101011010"; --    +226875    -262822
      WHEN 1197 => Ti := "000010111110001100110101000100011110001000010100"; --    +779061   +1171988
      WHEN 1198 => Ti := "000001000100101000101011111110011100111100000001"; --    +281131    -405759
      WHEN 1199 => Ti := "000000011110100000000010000011110001110111101110"; --    +124930    +990702
      WHEN 1200 => Ti := "000000101101111111101000111011010001100011111101"; --    +188392   -1238787
      WHEN 1201 => Ti := "000001000100100101011001111110010100111110010111"; --    +280921    -438377
      WHEN 1202 => Ti := "000001000001110001000110000001100111110110101011"; --    +269382    +425387
      WHEN 1203 => Ti := "111010101110110001101111111100000010111110111101"; --   -1381265   -1036355
      WHEN 1204 => Ti := "111011100111110110110110111101001011001111111011"; --   -1147466    -740357
      WHEN 1205 => Ti := "000010000011110110101111111111000101001111000000"; --    +540079    -240704
      WHEN 1206 => Ti := "111110001011100101010000000010110110001110000110"; --    -476848    +746374
      WHEN 1207 => Ti := "111111000011100000000111000000100111010001111001"; --    -247801    +160889
      WHEN 1208 => Ti := "000000011110000110100111000010111101101010111101"; --    +123303    +776893
      WHEN 1209 => Ti := "111111111111101000100000111101000010111000001001"; --      -1504    -774647
      WHEN 1210 => Ti := "111110100110000001010110000110001011101100111100"; --    -368554   +1620796
      WHEN 1211 => Ti := "111110111011010001011001000000011000111010011000"; --    -281511    +102040
      WHEN 1212 => Ti := "000001000011011011000011000001000101010000101011"; --    +276163    +283691
      WHEN 1213 => Ti := "000001000110011111010111111100100001000111111011"; --    +288727    -912901
      WHEN 1214 => Ti := "111100100111111101101000000000111100100111110011"; --    -884888    +248307
      WHEN 1215 => Ti := "000001101000111001111011111011001110001101011110"; --    +429691   -1252514
      WHEN 1216 => Ti := "000001100100010111000000000001010101110001110101"; --    +411072    +351349
      WHEN 1217 => Ti := "000011111000110100100111111110011100100111011101"; --   +1019175    -407075
      WHEN 1218 => Ti := "111100000100110110100101111101111011100110000011"; --   -1028699    -542333
      WHEN 1219 => Ti := "000100011101110110011011111110111010000111100001"; --   +1170843    -286239
      WHEN 1220 => Ti := "000000010101000111101000000000110000000110111011"; --     +86504    +197051
      WHEN 1221 => Ti := "111111001010101011010110111101001101001111010000"; --    -218410    -732208
      WHEN 1222 => Ti := "111101100011110110110000111110011101010010100001"; --    -639568    -404319
      WHEN 1223 => Ti := "111010101100011101001000000011001010001001101110"; --   -1390776    +828014
      WHEN 1224 => Ti := "000010010110001010100101111110100100000101110111"; --    +615077    -376457
      WHEN 1225 => Ti := "111111101100100111110111111111101000010010110100"; --     -79369     -97100
      WHEN 1226 => Ti := "000000000000011110001101000000000010100100111011"; --      +1933     +10555
      WHEN 1227 => Ti := "000001101111011110110111111010001010001000001110"; --    +456631   -1531378
      WHEN 1228 => Ti := "000001100111011100101011111111100010011111011011"; --    +423723    -120869
      WHEN 1229 => Ti := "111111111001001011001110111110111101101100001010"; --     -27954    -271606
      WHEN 1230 => Ti := "000001010001001010100000000011000101101110001110"; --    +332448    +809870
      WHEN 1231 => Ti := "000011011001110111000001111111000111000000000011"; --    +892353    -233469
      WHEN 1232 => Ti := "111110000001011001110001111111010010100000000010"; --    -518543    -186366
      WHEN 1233 => Ti := "111111011110110100001101111101010010110011110000"; --    -135923    -709392
      WHEN 1234 => Ti := "000010101111010101011111111101111010001010001010"; --    +718175    -548214
      WHEN 1235 => Ti := "000000001001010110111101000010100011110010011111"; --     +38333    +670879
      WHEN 1236 => Ti := "000001001101110100001011000011001010000101011010"; --    +318731    +827738
      WHEN 1237 => Ti := "111010100001110101100011111111110001010010011010"; --   -1434269     -60262
      WHEN 1238 => Ti := "000011100111011111100100111111010011010110010010"; --    +948196    -182894
      WHEN 1239 => Ti := "000011001001100001000100111110001111011100100111"; --    +825412    -461017
      WHEN 1240 => Ti := "000011100001111110110001000001000100011110001100"; --    +925617    +280460
      WHEN 1241 => Ti := "000001011011111110010001000010110011000000100011"; --    +376721    +733219
      WHEN 1242 => Ti := "111101101001001110111011000010111011110000100100"; --    -617541    +769060
      WHEN 1243 => Ti := "000000010000010100110001111101101000001011000001"; --     +66865    -621887
      WHEN 1244 => Ti := "000010110101001100110101000010100001010011010000"; --    +742197    +660688
      WHEN 1245 => Ti := "111111000010110100100101000000001111100101100100"; --    -250587     +63844
      WHEN 1246 => Ti := "000000101010110110001001000000001011111110111000"; --    +175497     +49080
      WHEN 1247 => Ti := "111110111000100010011001000001011101100111001001"; --    -292711    +383433
      WHEN 1248 => Ti := "000001010001001011010011000001101110111000110100"; --    +332499    +454196
      WHEN 1249 => Ti := "111101010111101001100000111011111100101001110110"; --    -689568   -1062282
      WHEN 1250 => Ti := "000001000101111101011100000100101101110111000100"; --    +286556   +1236420
      WHEN 1251 => Ti := "000001011001001010011111111101110111010110111001"; --    +365215    -559687
      WHEN 1252 => Ti := "000010101000010111000111111111100010100100110110"; --    +689607    -120522
      WHEN 1253 => Ti := "000001111111101101111001111010010010101100101010"; --    +523129   -1496278
      WHEN 1254 => Ti := "000101011001110111110011000000100011010110011011"; --   +1416691    +144795
      WHEN 1255 => Ti := "000000110110001101000011111111100101100110110010"; --    +222019    -108110
      WHEN 1256 => Ti := "000001000010100000111010000110011000011000111001"; --    +272442   +1672761
      WHEN 1257 => Ti := "111010011110100110000110111111110110000111000001"; --   -1447546     -40511
      WHEN 1258 => Ti := "000000001000110010101111110111000000011100011101"; --     +36015   -2357475
      WHEN 1259 => Ti := "000010010100110011011000000011001001111111010010"; --    +609496    +827346
      WHEN 1260 => Ti := "000010101110000101111010111110110111110011001100"; --    +713082    -295732
      WHEN 1261 => Ti := "000001011010010010111100000110110010001011100110"; --    +369852   +1778406
      WHEN 1262 => Ti := "000000110010001011101011000010000111011100001000"; --    +205547    +554760
      WHEN 1263 => Ti := "111011110110111100000101000010010111000011010111"; --   -1085691    +618711
      WHEN 1264 => Ti := "000101001110110000100101111011001100111001001100"; --   +1371173   -1257908
      WHEN 1265 => Ti := "111111110010100110110110000000001110111101110011"; --     -54858     +61299
      WHEN 1266 => Ti := "000000011000111000100110000010101111011100111111"; --    +101926    +718655
      WHEN 1267 => Ti := "111110101110100011100000000011110000110110011110"; --    -333600    +986526
      WHEN 1268 => Ti := "000011110111010101001011111110111001100000001100"; --   +1013067    -288756
      WHEN 1269 => Ti := "111010011111001010000111000010101100000010010000"; --   -1445241    +704656
      WHEN 1270 => Ti := "000000000110000010101101111011110111100011001011"; --     +24749   -1083189
      WHEN 1271 => Ti := "000011010000011100010101000010010100101100110010"; --    +853781    +609074
      WHEN 1272 => Ti := "111101100111001100010111000001101100000011101100"; --    -625897    +442604
      WHEN 1273 => Ti := "000000101010011001011101111111101100100101100111"; --    +173661     -79513
      WHEN 1274 => Ti := "000001101011010011101101111111100000000001110011"; --    +439533    -130957
      WHEN 1275 => Ti := "111111110100110110001111000001001010001111000010"; --     -45681    +304066
      WHEN 1276 => Ti := "111111010001111110110111111100111111101101001101"; --    -188489    -787635
      WHEN 1277 => Ti := "000000111000011001011010000001010101101101111001"; --    +231002    +351097
      WHEN 1278 => Ti := "000000011100001000010000111110100100101100100110"; --    +115216    -373978
      WHEN 1279 => Ti := "000010111011101011000101000010011101010110110010"; --    +768709    +644530
      WHEN 1280 => Ti := "000001011110101000010010111100011101111010111101"; --    +387602    -926019
      WHEN 1281 => Ti := "111111001100000110000000111101110101111110101110"; --    -212608    -565330
      WHEN 1282 => Ti := "111111011110011010011110000000010110010010100001"; --    -137570     +91297
      WHEN 1283 => Ti := "000001110100100100001100000011010100101101001111"; --    +477452    +871247
      WHEN 1284 => Ti := "111011110101101001111110000010011100010001100101"; --   -1090946    +640101
      WHEN 1285 => Ti := "000010101011100111101110111110010110011100101100"; --    +702958    -432340
      WHEN 1286 => Ti := "111111011100100100011101000000011010111011010001"; --    -145123    +110289
      WHEN 1287 => Ti := "111111011001101111101101111111000111111001000111"; --    -156691    -229817
      WHEN 1288 => Ti := "111111101011010101100000111110101001010001000001"; --     -84640    -355263
      WHEN 1289 => Ti := "000001010111100011001010111101101010100100001001"; --    +358602    -612087
      WHEN 1290 => Ti := "111100100100110110100100111110110010010001110010"; --    -897628    -318350
      WHEN 1291 => Ti := "000001010001110110111100111101111000010101101011"; --    +335292    -555669
      WHEN 1292 => Ti := "000011011110011000000101000010000000100011011101"; --    +910853    +526557
      WHEN 1293 => Ti := "111111100010101101001010111111001101010111100110"; --    -119990    -207386
      WHEN 1294 => Ti := "000000011101101011010011000011100110011101000110"; --    +121555    +943942
      WHEN 1295 => Ti := "000001101111000101010001000000001011100010111100"; --    +454993     +47292
      WHEN 1296 => Ti := "111001100100111100110111111100100101011000111011"; --   -1683657    -895429
      WHEN 1297 => Ti := "111111110100111100110110000000000110011111101001"; --     -45258     +26601
      WHEN 1298 => Ti := "000001110001111100011000000001100101000101000011"; --    +466712    +414019
      WHEN 1299 => Ti := "000000100101001000010001111100100110111110101001"; --    +152081    -888919
      WHEN 1300 => Ti := "111110001000111111010111000001100100001001110101"; --    -487465    +410229
      WHEN 1301 => Ti := "111111101000000000011110000010001000000011101010"; --     -98274    +557290
      WHEN 1302 => Ti := "111111110000101011001001111111101111101110101010"; --     -62775     -66646
      WHEN 1303 => Ti := "000101000010111100110110111111001001011011011110"; --   +1322806    -223522
      WHEN 1304 => Ti := "111101101100110111100011000101000000000111100111"; --    -602653   +1311207
      WHEN 1305 => Ti := "111110110101101000000010111111110000111000110010"; --    -304638     -61902
      WHEN 1306 => Ti := "111101000011000010001010111111100101000010010111"; --    -774006    -110441
      WHEN 1307 => Ti := "000100001000010101011000111010110000111001000100"; --   +1082712   -1372604
      WHEN 1308 => Ti := "111111011101000010111100111100011110111100010111"; --    -143172    -921833
      WHEN 1309 => Ti := "111111011110001100000001111011111000100100011111"; --    -138495   -1079009
      WHEN 1310 => Ti := "000000011000100001110001000000100100001011001110"; --    +100465    +148174
      WHEN 1311 => Ti := "111111111010111011010111111011100000000110111000"; --     -20777   -1179208
      WHEN 1312 => Ti := "000000101110000110101001111011101000011011010000"; --    +188841   -1145136
      WHEN 1313 => Ti := "111111101010001101001010000000001110011111010000"; --     -89270     +59344
      WHEN 1314 => Ti := "111110000111100000001011111010010111101010111010"; --    -493557   -1475910
      WHEN 1315 => Ti := "111101001010011011110110111010001100101111011101"; --    -743690   -1520675
      WHEN 1316 => Ti := "000000101010010000000111111111011111000100111110"; --    +173063    -134850
      WHEN 1317 => Ti := "000011101001011011010010111101000001110011110010"; --    +956114    -779022
      WHEN 1318 => Ti := "000000110011100001001001111010010010010010010001"; --    +211017   -1497967
      WHEN 1319 => Ti := "111110101100110110111010000001001100010110111000"; --    -340550    +312760
      WHEN 1320 => Ti := "111100110001100000011001111100010001011001101110"; --    -845799    -977298
      WHEN 1321 => Ti := "111110100100000010101110111110000111101101100001"; --    -376658    -492703
      WHEN 1322 => Ti := "000011000011001011010001000011101110101101101011"; --    +799441    +977771
      WHEN 1323 => Ti := "111110010111101011100110000010111001010100001010"; --    -427290    +759050
      WHEN 1324 => Ti := "111010011001111111100000000000110001100100011110"; --   -1466400    +203038
      WHEN 1325 => Ti := "111110111110001001100001000011101111010011001101"; --    -269727    +980173
      WHEN 1326 => Ti := "111101111011111100011010000010100011011100000110"; --    -540902    +669446
      WHEN 1327 => Ti := "111011110110010010110111000100000010110000111011"; --   -1088329   +1059899
      WHEN 1328 => Ti := "000001011100011010111110111100100110000011110100"; --    +378558    -892684
      WHEN 1329 => Ti := "000100000110000111110010111101110010110100011110"; --   +1073650    -578274
      WHEN 1330 => Ti := "111010011011101011100010111101000111010011110101"; --   -1459486    -756491
      WHEN 1331 => Ti := "111111110010011001011100000001101110111110110001"; --     -55716    +454577
      WHEN 1332 => Ti := "000100110100000100001111111011011111101101101111"; --   +1261839   -1180817
      WHEN 1333 => Ti := "111110000010001011101010000010100010111010011001"; --    -515350    +667289
      WHEN 1334 => Ti := "000001101110111011011111111011001010100101011111"; --    +454367   -1267361
      WHEN 1335 => Ti := "000000110010111010010110000001111010001010000111"; --    +208534    +500359
      WHEN 1336 => Ti := "000001010001010100100110111111001101100111001010"; --    +333094    -206390
      WHEN 1337 => Ti := "000000011000011010010101000000010000010100001110"; --     +99989     +66830
      WHEN 1338 => Ti := "000101000111101101010111111100001100010000001001"; --   +1342295    -998391
      WHEN 1339 => Ti := "111110101001110001010111111111010010010110100001"; --    -353193    -186975
      WHEN 1340 => Ti := "000001000001001010000000000000000010011111011010"; --    +266880     +10202
      WHEN 1341 => Ti := "111111001110110101011010111111111101011011011000"; --    -201382     -10536
      WHEN 1342 => Ti := "000001000011110110110111111011111001110110011001"; --    +277943   -1073767
      WHEN 1343 => Ti := "111011111001000111010110000110101010010100111101"; --   -1076778   +1746237
      WHEN 1344 => Ti := "000010001111001000010011000000100010011110100101"; --    +586259    +141221
      WHEN 1345 => Ti := "000000001101010001110101000000110011101100001110"; --     +54389    +211726
      WHEN 1346 => Ti := "000010111011001011110001111111011111011010111110"; --    +766705    -133442
      WHEN 1347 => Ti := "111110010010110010101110111111011110100010100101"; --    -447314    -137051
      WHEN 1348 => Ti := "000001111001100001010000111100100110111110001111"; --    +497744    -888945
      WHEN 1349 => Ti := "111110001110001011110000111011100100110101011110"; --    -466192   -1159842
      WHEN 1350 => Ti := "000000010011001101111111000001001010011010111101"; --     +78719    +304829
      WHEN 1351 => Ti := "000011111101110000100001111011100111100101101111"; --   +1039393   -1148561
      WHEN 1352 => Ti := "111111001100100100001100000100100101001101110011"; --    -210676   +1201011
      WHEN 1353 => Ti := "000001000000111000110010000010001010010100011110"; --    +265778    +566558
      WHEN 1354 => Ti := "000001001011001000110000000001110001101101010111"; --    +307760    +465751
      WHEN 1355 => Ti := "000010100000101010110111000101000111111101101101"; --    +658103   +1343341
      WHEN 1356 => Ti := "111101010111101111111110000000000000001110111000"; --    -689154       +952
      WHEN 1357 => Ti := "000101011010001111010100111100001110001101010010"; --   +1418196    -990382
      WHEN 1358 => Ti := "000001111110011011011010000001111001100101000110"; --    +517850    +497990
      WHEN 1359 => Ti := "111110011011111000110001000011000111010110001010"; --    -410063    +816522
      WHEN 1360 => Ti := "111100110101001100100011111110001001111001110100"; --    -830685    -483724
      WHEN 1361 => Ti := "000001111100100000111000000010111111110101001100"; --    +510008    +785740
      WHEN 1362 => Ti := "000010011111010100101100000010000101000101110010"; --    +652588    +545138
      WHEN 1363 => Ti := "111101000000101010110000000100101110011110000000"; --    -783696   +1238912
      WHEN 1364 => Ti := "000010010011111110000101111011101100000111110101"; --    +606085   -1129995
      WHEN 1365 => Ti := "111110111100001100011011000011001110100101000010"; --    -277733    +846146
      WHEN 1366 => Ti := "000011011111101100101111111101011010111111100011"; --    +916271    -675869
      WHEN 1367 => Ti := "000010001101100011011001111100010111000001010001"; --    +579801    -954287
      WHEN 1368 => Ti := "000001111000010101001101000000100111011010110000"; --    +492877    +161456
      WHEN 1369 => Ti := "000001011110011000111110111110000101111110001000"; --    +386622    -499832
      WHEN 1370 => Ti := "111111110001000110010000111110111000111111110000"; --     -61040    -290832
      WHEN 1371 => Ti := "000000011001001101100111000000110101101010110000"; --    +103271    +219824
      WHEN 1372 => Ti := "111010010000101100001110000001011100010000001001"; --   -1504498    +377865
      WHEN 1373 => Ti := "111100010111101001001101000011111011100011011010"; --    -951731   +1030362
      WHEN 1374 => Ti := "000001100111111100010100111111001010111011111110"; --    +425748    -217346
      WHEN 1375 => Ti := "000001110100111111100010000110010111000010111010"; --    +479202   +1667258
      WHEN 1376 => Ti := "000010100111011110010000000010110000100111110010"; --    +685968    +723442
      WHEN 1377 => Ti := "000010001100010110111101111101101110100000110111"; --    +574909    -595913
      WHEN 1378 => Ti := "111110001101010111111111111111111000111100101100"; --    -469505     -28884
      WHEN 1379 => Ti := "000000001111101111100101111111001001011111010011"; --     +64485    -223277
      WHEN 1380 => Ti := "000001010000001011000100111111100010111001110111"; --    +328388    -119177
      WHEN 1381 => Ti := "000001011101100101100011111100011110010010111010"; --    +383331    -924486
      WHEN 1382 => Ti := "000011100100001000101101111110011100001111101101"; --    +934445    -408595
      WHEN 1383 => Ti := "111110111001001010101100111110101100011111111110"; --    -290132    -342018
      WHEN 1384 => Ti := "000000110011001111110010111011011110000110110011"; --    +209906   -1187405
      WHEN 1385 => Ti := "111110011000101100011011111101010010011011001100"; --    -423141    -710964
      WHEN 1386 => Ti := "000000100111101101101001111111100100101100101001"; --    +162665    -111831
      WHEN 1387 => Ti := "111100111001110000101101000011101111000100001001"; --    -811987    +979209
      WHEN 1388 => Ti := "111111010101001111110111000010010101010101111101"; --    -175113    +611709
      WHEN 1389 => Ti := "000010101010110100010110000001000010011100111101"; --    +699670    +272189
      WHEN 1390 => Ti := "000010110010011101001101000001100010101010100001"; --    +730957    +404129
      WHEN 1391 => Ti := "000000011101000100100000111110101110010100100010"; --    +119072    -334558
      WHEN 1392 => Ti := "111100110110111100111100111101010001011000110011"; --    -823492    -715213
      WHEN 1393 => Ti := "000000111000101001001101111111010101101110010101"; --    +232013    -173163
      WHEN 1394 => Ti := "111110001011001100011011111100101011011110100110"; --    -478437    -870490
      WHEN 1395 => Ti := "000100011001000001100001111101000010111100100001"; --   +1151073    -774367
      WHEN 1396 => Ti := "000001010111101101100111111111101000110101011011"; --    +359271     -94885
      WHEN 1397 => Ti := "111110100000001101101101111110010101011000100101"; --    -392339    -436699
      WHEN 1398 => Ti := "000110011110001011111100111110100001001010000001"; --   +1696508    -388479
      WHEN 1399 => Ti := "000011101100000100101010000101110110101001110100"; --    +966954   +1534580
      WHEN 1400 => Ti := "000001101111101110101010111101001011000110000101"; --    +457642    -740987
      WHEN 1401 => Ti := "111110000000101100010100000011110111100011101110"; --    -521452   +1013998
      WHEN 1402 => Ti := "000000010000010010001101000011011100110011111010"; --     +66701    +904442
      WHEN 1403 => Ti := "111111010101110000100100000000001101100100111101"; --    -173020     +55613
      WHEN 1404 => Ti := "000010000101001100010100000010010010100111100100"; --    +545556    +600548
      WHEN 1405 => Ti := "111111110000011000101100000010100110100011001100"; --     -63956    +682188
      WHEN 1406 => Ti := "111110100101011001100111111101101011100001101010"; --    -371097    -608150
      WHEN 1407 => Ti := "000011011010111000000111111111011101111011011011"; --    +896519    -139557
      WHEN 1408 => Ti := "111100101000111001011011111100100110100100101101"; --    -881061    -890579
      WHEN 1409 => Ti := "000010010101001001000110111110100011001010000110"; --    +610886    -380282
      WHEN 1410 => Ti := "111111010011010010110000000001001101010011011101"; --    -183120    +316637
      WHEN 1411 => Ti := "000001010111011111101101111111101001101011001100"; --    +358381     -91444
      WHEN 1412 => Ti := "000100110110001010100000000000000011101100001011"; --   +1270432     +15115
      WHEN 1413 => Ti := "111111100110110101110010111011111111101110101001"; --    -103054   -1049687
      WHEN 1414 => Ti := "111111111000111110001101000000000000001101111111"; --     -28787       +895
      WHEN 1415 => Ti := "111110110111011110101111000010000101101001000110"; --    -297041    +547398
      WHEN 1416 => Ti := "000010001001001111100000000001100010110101110000"; --    +562144    +404848
      WHEN 1417 => Ti := "000100111000111101010000000010000011101001011010"; --   +1281872    +539226
      WHEN 1418 => Ti := "000101001011110000000010000000101111001001010011"; --   +1358850    +193107
      WHEN 1419 => Ti := "111110111101111100111111000001010110111110011000"; --    -270529    +356248
      WHEN 1420 => Ti := "111100011010111011011001000000000011110101000001"; --    -938279     +15681
      WHEN 1421 => Ti := "111101100111001001000011111110111100001100011010"; --    -626109    -277734
      WHEN 1422 => Ti := "000010000010111110111001000000000000110111011000"; --    +536505      +3544
      WHEN 1423 => Ti := "000001111101111101000111111101011011010110111101"; --    +515911    -674371
      WHEN 1424 => Ti := "000000101010100010101100111011100100010001010011"; --    +174252   -1162157
      WHEN 1425 => Ti := "111011111011110100001001000000100001011010100101"; --   -1065719    +136869
      WHEN 1426 => Ti := "111111011001110000100111000000110111100001110010"; --    -156633    +227442
      WHEN 1427 => Ti := "111100101011001000001010000010111010001000011100"; --    -871926    +762396
      WHEN 1428 => Ti := "111111011000011110001010111100111110010001110100"; --    -161910    -793484
      WHEN 1429 => Ti := "111111110010110110010010000000011110000011010011"; --     -53870    +123091
      WHEN 1430 => Ti := "111111000010111101001010111111011100011101011101"; --    -250038    -145571
      WHEN 1431 => Ti := "111100010110100010011010111100011010101110111010"; --    -956262    -939078
      WHEN 1432 => Ti := "111101100100111000101011000001011010011110101111"; --    -635349    +370607
      WHEN 1433 => Ti := "111100101110110111001011000000001100111101101110"; --    -856629     +53102
      WHEN 1434 => Ti := "111101001010011110001111111100100110110111100110"; --    -743537    -889370
      WHEN 1435 => Ti := "000000011000011010010101000011010010110110110010"; --     +99989    +863666
      WHEN 1436 => Ti := "111011010110111001100100000010100001101011010011"; --   -1216924    +662227
      WHEN 1437 => Ti := "000101000000101000000010000001111110101010111111"; --   +1313282    +518847
      WHEN 1438 => Ti := "111101101101001101000111111011110111010011111100"; --    -601273   -1084164
      WHEN 1439 => Ti := "111110101111000011101000111101100001011001001101"; --    -331544    -649651
      WHEN 1440 => Ti := "111111111010001101000011000001100000100010000001"; --     -23741    +395393
      WHEN 1441 => Ti := "111101100101010000110000000101100001111101100110"; --    -633808   +1449830
      WHEN 1442 => Ti := "111110111010101110111110111010011011100100100101"; --    -283714   -1459931
      WHEN 1443 => Ti := "000101000011001111000100000001010101100010011010"; --   +1323972    +350362
      WHEN 1444 => Ti := "000010000011101111101110111011001100111101100111"; --    +539630   -1257625
      WHEN 1445 => Ti := "000001001011110001010110111111010010100111101101"; --    +310358    -185875
      WHEN 1446 => Ti := "000000010011101000100101000010011100000001011001"; --     +80421    +639065
      WHEN 1447 => Ti := "000101100101101000101110000001100100001001010110"; --   +1464878    +410198
      WHEN 1448 => Ti := "000110011111110100100111000010100001100110000111"; --   +1703207    +661895
      WHEN 1449 => Ti := "111110110010001100001010111101111100101100001001"; --    -318710    -537847
      WHEN 1450 => Ti := "000000010000101010111100000010100000110111011011"; --     +68284    +658907
      WHEN 1451 => Ti := "000100010011101111011111000001000100100110011100"; --   +1129439    +280988
      WHEN 1452 => Ti := "000011001011001101001111000000011000111000010010"; --    +832335    +101906
      WHEN 1453 => Ti := "111111011000010101101000111110110100111010111111"; --    -162456    -307521
      WHEN 1454 => Ti := "111111001100000001000000000001000100101111010110"; --    -212928    +281558
      WHEN 1455 => Ti := "111110100100101100000010000001110010111100001110"; --    -374014    +470798
      WHEN 1456 => Ti := "000011010010001001001010111110100011011110101010"; --    +860746    -378966
      WHEN 1457 => Ti := "111010100111000100110100000000010110010111110100"; --   -1412812     +91636
      WHEN 1458 => Ti := "111110010111110110100100000001011010110110101111"; --    -426588    +372143
      WHEN 1459 => Ti := "000000011011100010110001111111011100111101011111"; --    +112817    -143521
      WHEN 1460 => Ti := "000001011000100010111101111100001001110011100111"; --    +362685   -1008409
      WHEN 1461 => Ti := "111101111110101110110101000100101101000101100001"; --    -529483   +1233249
      WHEN 1462 => Ti := "000100000101111001100100000001000100011000100010"; --   +1072740    +280098
      WHEN 1463 => Ti := "111101000010101010010001000010101010001101111011"; --    -775535    +697211
      WHEN 1464 => Ti := "000010110010111000001101111100001111000100001011"; --    +732685    -986869
      WHEN 1465 => Ti := "111111100101110110011010111110100111010100010100"; --    -107110    -363244
      WHEN 1466 => Ti := "111011010001110111011010111110110100100001010101"; --   -1237542    -309163
      WHEN 1467 => Ti := "111110010010100111100110111101010111010010110111"; --    -448026    -691017
      WHEN 1468 => Ti := "000000011010101110011111111111110001111111010110"; --    +109471     -57386
      WHEN 1469 => Ti := "000100011001011010000011111110000011001100010100"; --   +1152643    -511212
      WHEN 1470 => Ti := "000000101001100010100110000011000111010010100001"; --    +170150    +816289
      WHEN 1471 => Ti := "111101011101001110100010111111001000100011001100"; --    -666718    -227124
      WHEN 1472 => Ti := "000001010100110011000100000011001011000000110011"; --    +347332    +831539
      WHEN 1473 => Ti := "000011011101100100011001000000010000010011111010"; --    +907545     +66810
      WHEN 1474 => Ti := "111110000110001110111001000001110001100001110001"; --    -498759    +465009
      WHEN 1475 => Ti := "000000010110010110000001111111100000100110101100"; --     +91521    -128596
      WHEN 1476 => Ti := "111011000101100110010100111110111100001010100011"; --   -1287788    -277853
      WHEN 1477 => Ti := "000011001101101101010001000100100110000011001011"; --    +842577   +1204427
      WHEN 1478 => Ti := "111101111101101100011101111110100001101100100011"; --    -533731    -386269
      WHEN 1479 => Ti := "111100111010000010000110000000110010110110100110"; --    -810874    +208294
      WHEN 1480 => Ti := "000000000010010101000101111000111110101001110110"; --      +9541   -1840522
      WHEN 1481 => Ti := "000000101110010010100011111110010001011010100000"; --    +189603    -452960
      WHEN 1482 => Ti := "111111101100111100111001000000110010101100001010"; --     -78023    +207626
      WHEN 1483 => Ti := "111110001100110000100110111111101101001100101010"; --    -472026     -77014
      WHEN 1484 => Ti := "111001111101111111000010111001000110101000011111"; --   -1581118   -1807841
      WHEN 1485 => Ti := "000010110000111101011000000000000100011100100111"; --    +724824     +18215
      WHEN 1486 => Ti := "111101111011011001011011111111110101000111001111"; --    -543141     -44593
      WHEN 1487 => Ti := "000100111000011100100110111101110001111001110011"; --   +1279782    -582029
      WHEN 1488 => Ti := "111111001011111111010111111110101100111000011011"; --    -213033    -340453
      WHEN 1489 => Ti := "111101100001001100110111000001110111001011111101"; --    -650441    +488189
      WHEN 1490 => Ti := "000000011001001000000001111110110000100000011011"; --    +102913    -325605
      WHEN 1491 => Ti := "000000000000110110011011000001111010100000011001"; --      +3483    +501785
      WHEN 1492 => Ti := "000001010010111100100001000101001010110010001100"; --    +339745   +1354892
      WHEN 1493 => Ti := "000101100000101000001000111101010000111010010001"; --   +1444360    -717167
      WHEN 1494 => Ti := "111110000000011010101011111101100011011100101101"; --    -522581    -641235
      WHEN 1495 => Ti := "000101000100111001000011000001000001101001110001"; --   +1330755    +268913
      WHEN 1496 => Ti := "000001111011110100111010000011110100100011101100"; --    +507194   +1001708
      WHEN 1497 => Ti := "111111101100110111000010000000111110100011110010"; --     -78398    +256242
      WHEN 1498 => Ti := "111100010010110100100100111111010111111110101010"; --    -971484    -163926
      WHEN 1499 => Ti := "111011011001111100101010000000011000001101110110"; --   -1204438     +99190
      WHEN 1500 => Ti := "111111111110010110000100111111110000101101111000"; --      -6780     -62600
      WHEN 1501 => Ti := "111101010001110011110001111111000010100010011111"; --    -713487    -251745
      WHEN 1502 => Ti := "111100110011101110010000000011101010000101111001"; --    -836720    +958841
      WHEN 1503 => Ti := "000001010111000011110001111110001100101110011111"; --    +356593    -472161
      WHEN 1504 => Ti := "000000101110111010101111111101101110111001000111"; --    +192175    -594361
      WHEN 1505 => Ti := "000110110011100010101011000001010001110011100011"; --   +1783979    +335075
      WHEN 1506 => Ti := "111011100010010110111110111101100110000011101001"; --   -1169986    -630551
      WHEN 1507 => Ti := "111111111011111000111101000000001000000010010011"; --     -16835     +32915
      WHEN 1508 => Ti := "000000011010101010100001111111110111101101011101"; --    +109217     -33955
      WHEN 1509 => Ti := "111111011110101100001100111110001100010111100111"; --    -136436    -473625
      WHEN 1510 => Ti := "000100000101101101110111111011010000100010100001"; --   +1071991   -1242975
      WHEN 1511 => Ti := "111101001100011000011100000011010011111111010110"; --    -735716    +868310
      WHEN 1512 => Ti := "000011000111001111000110111110100011110111011001"; --    +816070    -377383
      WHEN 1513 => Ti := "111110010110010111111111000000100000100111010000"; --    -432641    +133584
      WHEN 1514 => Ti := "111100110000101100110001111101100001010111000010"; --    -849103    -649790
      WHEN 1515 => Ti := "000001100100001010000001111010011011101110001111"; --    +410241   -1459313
      WHEN 1516 => Ti := "000000001010000101000101110111111000001100010000"; --     +41285   -2129136
      WHEN 1517 => Ti := "111111001011111100000111111101000110010010101000"; --    -213241    -760664
      WHEN 1518 => Ti := "111100110111010000110111000010001010011111111000"; --    -822217    +567288
      WHEN 1519 => Ti := "000000011000111000100000111110111111000110010110"; --    +101920    -265834
      WHEN 1520 => Ti := "111110110011110010101110111111011111010111110001"; --    -312146    -133647
      WHEN 1521 => Ti := "000001000001110110000111111101000101011111001000"; --    +269703    -763960
      WHEN 1522 => Ti := "111010100000100000011001111111010100001000010111"; --   -1439719    -179689
      WHEN 1523 => Ti := "111101100101110101100110000011000010111000100011"; --    -631450    +798243
      WHEN 1524 => Ti := "111110001000001111001100000100011101000100101000"; --    -490548   +1167656
      WHEN 1525 => Ti := "111101101010101011001101111100110000110111000011"; --    -611635    -848445
      WHEN 1526 => Ti := "111011100010100100010001111100111010110101111110"; --   -1169135    -807554
      WHEN 1527 => Ti := "111101010000010111111110111101000111111001111011"; --    -719362    -754053
      WHEN 1528 => Ti := "000001011010001011101110111100100111111001001000"; --    +369390    -885176
      WHEN 1529 => Ti := "000000110000100011111011000000000000010010111001"; --    +198907      +1209
      WHEN 1530 => Ti := "000001011111001100000000000001101100110001000100"; --    +389888    +445508
      WHEN 1531 => Ti := "111111010110110101100101111110011111011110111111"; --    -168603    -395329
      WHEN 1532 => Ti := "000010001000000000011100111100000111111011001100"; --    +557084   -1016116
      WHEN 1533 => Ti := "000001100001110110100111111111110111110111101110"; --    +400807     -33298
      WHEN 1534 => Ti := "000001110011000001001111111100101101101000000010"; --    +471119    -861694
      WHEN 1535 => Ti := "111110011010011101101110111100110000010010010010"; --    -415890    -850798
      WHEN 1536 => Ti := "000000100011110100111101000001110100000110011000"; --    +146749    +475544
      WHEN 1537 => Ti := "111110010000100110100110111100010111100101110110"; --    -456282    -951946
      WHEN 1538 => Ti := "111111101010100101001000000010101000111100111111"; --     -87736    +692031
      WHEN 1539 => Ti := "000000110101001000010011000000111101001111101100"; --    +217619    +250860
      WHEN 1540 => Ti := "111110011010001100101111111101100001001001110100"; --    -416977    -650636
      WHEN 1541 => Ti := "111111010001100110110111000000100111111001100001"; --    -190025    +163425
      WHEN 1542 => Ti := "111111001100001111110111111001011110101101111000"; --    -211977   -1709192
      WHEN 1543 => Ti := "000000111101110001100110111110000110100111000111"; --    +253030    -497209
      WHEN 1544 => Ti := "000011111001010000100000111101100001100100111111"; --   +1020960    -648897
      WHEN 1545 => Ti := "111110101100110100010000000000101100001101000001"; --    -340720    +181057
      WHEN 1546 => Ti := "111110001110000111101100000010000001011000110001"; --    -466452    +529969
      WHEN 1547 => Ti := "111110110011100110111000111111001100000100110001"; --    -312904    -212687
      WHEN 1548 => Ti := "111111100011000010110000111101111110101011110111"; --    -118608    -529673
      WHEN 1549 => Ti := "111101101010010111110111000000011101101011110111"; --    -612873    +121591
      WHEN 1550 => Ti := "111110110001000100011000111111100001011010000100"; --    -323304    -125308
      WHEN 1551 => Ti := "000000001111010101000111111001000101111111111001"; --     +62791   -1810439
      WHEN 1552 => Ti := "111110000111101000111100111011111001010100001111"; --    -492996   -1075953
      WHEN 1553 => Ti := "000010101001001011001100000000110001101011101101"; --    +692940    +203501
      WHEN 1554 => Ti := "111111110100010111111010111111010110000100110101"; --     -47622    -171723
      WHEN 1555 => Ti := "111111001100100100010010000010010010001010000010"; --    -210670    +598658
      WHEN 1556 => Ti := "000000000000010101101110111011010010110010001101"; --      +1390   -1233779
      WHEN 1557 => Ti := "000010101111010111101100000001110100110000101100"; --    +718316    +478252
      WHEN 1558 => Ti := "000000001100101001001110000010001111001010111110"; --     +51790    +586430
      WHEN 1559 => Ti := "000000110100100010100101111110000100110100110010"; --    +215205    -504526
      WHEN 1560 => Ti := "000000100010011110010010000010111111100100011101"; --    +141202    +784669
      WHEN 1561 => Ti := "000100011101101100010011111110100010011110000110"; --   +1170195    -383098
      WHEN 1562 => Ti := "000000000110100011000100111111101100000100000010"; --     +26820     -81662
      WHEN 1563 => Ti := "111111100011100101101100111110001111011110100110"; --    -116372    -460890
      WHEN 1564 => Ti := "000000101110010011111010000010011010101001101000"; --    +189690    +633448
      WHEN 1565 => Ti := "000001111111110010110110000000000100010111100000"; --    +523446     +17888
      WHEN 1566 => Ti := "000010001000111110011001111100000001110100101001"; --    +561049   -1041111
      WHEN 1567 => Ti := "111110000001111111000011000010011000101101110111"; --    -516157    +625527
      WHEN 1568 => Ti := "111100110111010110011100111111010010000101000110"; --    -821860    -188090
      WHEN 1569 => Ti := "111111100111000010101100111101100111011001101111"; --    -102228    -625041
      WHEN 1570 => Ti := "111110101111101100110000000001110110101000000100"; --    -328912    +485892
      WHEN 1571 => Ti := "000001110010011000010100111111100011000011101100"; --    +468500    -118548
      WHEN 1572 => Ti := "000010110000010001011111111111101011101110011110"; --    +722015     -83042
      WHEN 1573 => Ti := "111111101011001011100110111111001000011110000010"; --     -85274    -227454
      WHEN 1574 => Ti := "111011110101001101010110000001101110100010111111"; --   -1092778    +452799
      WHEN 1575 => Ti := "000001101001001110010000000011001101110011101111"; --    +430992    +842991
      WHEN 1576 => Ti := "111101010110000101011111111101000001110111100101"; --    -695969    -778779
      WHEN 1577 => Ti := "000001010000101101010111111111100111110101000110"; --    +330583     -99002
      WHEN 1578 => Ti := "000000111010010111111000111110000101110011010000"; --    +239096    -500528
      WHEN 1579 => Ti := "111101000001100101001000000001100010000010111010"; --    -779960    +401594
      WHEN 1580 => Ti := "000001101011101101001010111101101100010001110101"; --    +441162    -605067
      WHEN 1581 => Ti := "000000000011001000110101001000110111011011110000"; --     +12853   +2324208
      WHEN 1582 => Ti := "111110100111101101101100000010010001011100100100"; --    -361620    +595748
      WHEN 1583 => Ti := "000011110101101000101110000001001010011011110011"; --   +1006126    +304883
      WHEN 1584 => Ti := "000001010111000100000011000001010101110100100010"; --    +356611    +351522
      WHEN 1585 => Ti := "000010110010110111001111111100001110001011000000"; --    +732623    -990528
      WHEN 1586 => Ti := "111111110001101110111101111101110010110101110111"; --     -58435    -578185
      WHEN 1587 => Ti := "111111011000001110001101000000111110001000110110"; --    -162931    +254518
      WHEN 1588 => Ti := "111111010000110000001110111111101011111000110100"; --    -193522     -82380
      WHEN 1589 => Ti := "000000000001111101110110111011001101011110101000"; --      +8054   -1255512
      WHEN 1590 => Ti := "111111100001101001000110111110011001010100101010"; --    -124346    -420566
      WHEN 1591 => Ti := "111110000111000111010101111111011100010110011001"; --    -495147    -146023
      WHEN 1592 => Ti := "000000101001001000000111000011101010001010101101"; --    +168455    +959149
      WHEN 1593 => Ti := "111110111110010101110110111011001010100011000001"; --    -268938   -1267519
      WHEN 1594 => Ti := "000000110111000100111111111111101000000010100001"; --    +225599     -98143
      WHEN 1595 => Ti := "000001011011111000101011000001101101011000011010"; --    +376363    +448026
      WHEN 1596 => Ti := "111110101000100011011011111101111001011010110101"; --    -358181    -551243
      WHEN 1597 => Ti := "000010110111010110001111000000001101111011101111"; --    +750991     +57071
      WHEN 1598 => Ti := "111111101001100010001101000011011110010111000010"; --     -92019    +910786
      WHEN 1599 => Ti := "000000000000100011001001000011100100111100100011"; --      +2249    +937763
      WHEN 1600 => Ti := "000001011101100000000110111010011110101011011011"; --    +382982   -1447205
      WHEN 1601 => Ti := "111101111101111000011000111100100110100101000111"; --    -532968    -890553
      WHEN 1602 => Ti := "111011011011111110001011000000011111000101010011"; --   -1196149    +127315
      WHEN 1603 => Ti := "111011011111010001001011000100010110110001100101"; --   -1182645   +1141861
      WHEN 1604 => Ti := "000000010010001110000001000010100001010110111110"; --     +74625    +660926
      WHEN 1605 => Ti := "000011101111100100010111000000100110100100111100"; --    +981271    +158012
      WHEN 1606 => Ti := "000000000010001110011001000010011111110000010001"; --      +9113    +654353
      WHEN 1607 => Ti := "000100111001110001001100111111011110001011100110"; --   +1285196    -138522
      WHEN 1608 => Ti := "000000110110111101011000111100111010001110001110"; --    +225112    -810098
      WHEN 1609 => Ti := "111110011011001011110111000010000101100000001101"; --    -412937    +546829
      WHEN 1610 => Ti := "000101001111100111010110000001000101010101100101"; --   +1374678    +284005
      WHEN 1611 => Ti := "111111010110010011010101111110001000010111110000"; --    -170795    -490000
      WHEN 1612 => Ti := "111110011101101100010111111111111101010001001010"; --    -402665     -11190
      WHEN 1613 => Ti := "000010111111110100000110000001011110101101111101"; --    +785670    +387965
      WHEN 1614 => Ti := "111110000000010000111101000100101000101001100000"; --    -523203   +1215072
      WHEN 1615 => Ti := "111111001011010101010101111011010000011000011000"; --    -215723   -1243624
      WHEN 1616 => Ti := "000011011101001101110010111101110000010101111001"; --    +906098    -588423
      WHEN 1617 => Ti := "111100001111110101010010111111110100111110011011"; --    -983726     -45157
      WHEN 1618 => Ti := "000000011111001110001101000000011111010010101010"; --    +127885    +128170
      WHEN 1619 => Ti := "111111011001000110001110111100000111100010111110"; --    -159346   -1017666
      WHEN 1620 => Ti := "000001001001000001001101000000111110110100001100"; --    +299085    +257292
      WHEN 1621 => Ti := "111101011010000010101100111101101111011101000100"; --    -679764    -592060
      WHEN 1622 => Ti := "111101000111101001101111000001001000011011100001"; --    -755089    +296673
      WHEN 1623 => Ti := "000001100001110101000110111111100000001011001000"; --    +400710    -130360
      WHEN 1624 => Ti := "000100110000011011001101000000010111110111100011"; --   +1246925     +97763
      WHEN 1625 => Ti := "111101100100011000101100111101001110011000010000"; --    -637396    -727536
      WHEN 1626 => Ti := "000010101110000001011101000000010111001011101011"; --    +712797     +94955
      WHEN 1627 => Ti := "111110010110111111010011000010100001010101101001"; --    -430125    +660841
      WHEN 1628 => Ti := "111111000011000011001011000000010100000010110100"; --    -249653     +82100
      WHEN 1629 => Ti := "111111000110010001101010000011101101100111111111"; --    -236438    +973311
      WHEN 1630 => Ti := "111110111111001000100010000100101000011111111100"; --    -265694   +1214460
      WHEN 1631 => Ti := "111100011100101000110110000001011111100011000010"; --    -931274    +391362
      WHEN 1632 => Ti := "000010010110100011001001000010110011100110011110"; --    +616649    +735646
      WHEN 1633 => Ti := "000001111001011011000010111111010110000100001111"; --    +497346    -171761
      WHEN 1634 => Ti := "000100001110100111101000000000010110111000001100"; --   +1108456     +93708
      WHEN 1635 => Ti := "111111000000111101100010111001110001111010001110"; --    -258206   -1630578
      WHEN 1636 => Ti := "000000110000000000001011111100100110101010011111"; --    +196619    -890209
      WHEN 1637 => Ti := "000101011010000100000001000000010011100111000100"; --   +1417473     +80324
      WHEN 1638 => Ti := "111111111011111010011111111111000101100110010010"; --     -16737    -239214
      WHEN 1639 => Ti := "000001101011111010011001000010011111010111000111"; --    +442009    +652743
      WHEN 1640 => Ti := "111101111110011101101101000001001100101001111011"; --    -530579    +313979
      WHEN 1641 => Ti := "111100111110001100101001000001001110111011100011"; --    -793815    +323299
      WHEN 1642 => Ti := "000010010011110000101010000011000101010100001110"; --    +605226    +808206
      WHEN 1643 => Ti := "111100001111110100111110111100101101111110000000"; --    -983746    -860288
      WHEN 1644 => Ti := "000000010011001111011111111110011111110101011101"; --     +78815    -393891
      WHEN 1645 => Ti := "000001111101110101000101111010110010001101101001"; --    +515397   -1367191
      WHEN 1646 => Ti := "000000001111100111001101000000101111011011100101"; --     +63949    +194277
      WHEN 1647 => Ti := "111101001000101001000101000011010111110111001000"; --    -751035    +884168
      WHEN 1648 => Ti := "000001100001001011001010000010110010100000001100"; --    +398026    +731148
      WHEN 1649 => Ti := "000010101010110100000100000100001111010100011001"; --    +699652   +1111321
      WHEN 1650 => Ti := "111101010011010110011100000001011000000101000000"; --    -707172    +360768
      WHEN 1651 => Ti := "111110110011011101111100000000001001110100011000"; --    -313476     +40216
      WHEN 1652 => Ti := "111110010001100100110111000000100011000010111111"; --    -452297    +143551
      WHEN 1653 => Ti := "000001001010100101011010000010001111110100101010"; --    +305498    +589098
      WHEN 1654 => Ti := "111111101100110010010111000011100110011010000010"; --     -78697    +943746
      WHEN 1655 => Ti := "000001001011001001011111000010011010011011010010"; --    +307807    +632530
      WHEN 1656 => Ti := "111010111011010011011111000001000000111101010101"; --   -1329953    +266069
      WHEN 1657 => Ti := "111101010000010010000011000000001011111110011110"; --    -719741     +49054
      WHEN 1658 => Ti := "000101001011100110100110000001001100010011001100"; --   +1358246    +312524
      WHEN 1659 => Ti := "111110110001010000011011000010001001101100011011"; --    -322533    +563995
      WHEN 1660 => Ti := "000000010001000011000011111101101000000100100010"; --     +69827    -622302
      WHEN 1661 => Ti := "111101111111110111111100111111001011110111001010"; --    -524804    -213558
      WHEN 1662 => Ti := "111111000111011110000101000000010110010010001010"; --    -231547     +91274
      WHEN 1663 => Ti := "111111111011111101000010000010000001011100011010"; --     -16574    +530202
      WHEN 1664 => Ti := "111111111110011001001101000000000110111110111011"; --      -6579     +28603
      WHEN 1665 => Ti := "000000101010011111011011111010111111001000011010"; --    +174043   -1314278
      WHEN 1666 => Ti := "000001000101110001101011111111111101000100100010"; --    +285803     -11998
      WHEN 1667 => Ti := "000000110111011001110110111010110101111110011100"; --    +226934   -1351780
      WHEN 1668 => Ti := "111010111100001101000110000010110010110101101110"; --   -1326266    +732526
      WHEN 1669 => Ti := "111100111000101010100001000010000011010001000110"; --    -816479    +537670
      WHEN 1670 => Ti := "000000010110000000001101000011011101010101101100"; --     +90125    +906604
      WHEN 1671 => Ti := "000001100101100110100101111110001011100110001000"; --    +416165    -476792
      WHEN 1672 => Ti := "111101101110011001111100000011100001101011010101"; --    -596356    +924373
      WHEN 1673 => Ti := "000010011101001101100111000101010111110100001101"; --    +643943   +1408269
      WHEN 1674 => Ti := "000001001101111100100010111011000101101110010000"; --    +319266   -1287280
      WHEN 1675 => Ti := "000010101110100011111101111110001001110000000101"; --    +715005    -484347
      WHEN 1676 => Ti := "000000110110000000000111000000100001010101100110"; --    +221191    +136550
      WHEN 1677 => Ti := "000000010010110010000001000000011111111000001101"; --     +76929    +130573
      WHEN 1678 => Ti := "000010100100011110101010111110100000001011010010"; --    +673706    -392494
      WHEN 1679 => Ti := "000011001011010011001001000010101111011110101010"; --    +832713    +718762
      WHEN 1680 => Ti := "111111011101011010110011000001011010101011110100"; --    -141645    +371444
      WHEN 1681 => Ti := "111101000011111000100000111101110011010100000011"; --    -770528    -576253
      WHEN 1682 => Ti := "111111001111100010000110111010101010000000010010"; --    -198522   -1400814
      WHEN 1683 => Ti := "000110111000101100101111000001111100000010010010"; --   +1805103    +508050
      WHEN 1684 => Ti := "000110101100101010010011000000011101110001011100"; --   +1755795    +121948
      WHEN 1685 => Ti := "111011011111111101111011000000001011110000000010"; --   -1179781     +48130
      WHEN 1686 => Ti := "000010111010001011000110111111111000111101110100"; --    +762566     -28812
      WHEN 1687 => Ti := "111111010110000111111110111101010011100101101010"; --    -171522    -706198
      WHEN 1688 => Ti := "000000001001110101101000000001101100101011100011"; --     +40296    +445155
      WHEN 1689 => Ti := "000000001110011111010101111101010110100000001001"; --     +59349    -694263
      WHEN 1690 => Ti := "111101110100101011110010000100001001110100011111"; --    -570638   +1088799
      WHEN 1691 => Ti := "000011110010010001110010000001001110000000000100"; --    +992370    +319492
      WHEN 1692 => Ti := "000001100110100000100011111101100110001111011010"; --    +419875    -629798
      WHEN 1693 => Ti := "111100110011010000110110111101111110010000110111"; --    -838602    -531401
      WHEN 1694 => Ti := "000001000110101011100000111111000111100101001001"; --    +289504    -231095
      WHEN 1695 => Ti := "000000101101110110001011000001000111000010101100"; --    +187787    +290988
      WHEN 1696 => Ti := "000000011010111000111001000001011010101100001001"; --    +110137    +371465
      WHEN 1697 => Ti := "111110000000101110110101111111001001110011101111"; --    -521291    -221969
      WHEN 1698 => Ti := "111111010011000111101101111011110111100000010010"; --    -183827   -1083374
      WHEN 1699 => Ti := "111100000010110010110001000010110001011101111000"; --   -1037135    +726904
      WHEN 1700 => Ti := "111111000001100110101000000100010000010100000011"; --    -255576   +1115395
      WHEN 1701 => Ti := "000000011000000101011000000000100000101001110100"; --     +98648    +133748
      WHEN 1702 => Ti := "111111100000001100010010111100001011001010010001"; --    -130286   -1002863
      WHEN 1703 => Ti := "111110110011110000000010111111001110011110111111"; --    -312318    -202817
      WHEN 1704 => Ti := "000000100101001110010011111101000110100101111001"; --    +152467    -759431
      WHEN 1705 => Ti := "111101100111011110111011000000000001100100000101"; --    -624709      +6405
      WHEN 1706 => Ti := "111100010010101110110010111011101100011111001111"; --    -971854   -1128497
      WHEN 1707 => Ti := "111111100110011101101100000001101110001111011111"; --    -104596    +451551
      WHEN 1708 => Ti := "111111111010111110010111111110110000000010000100"; --     -20585    -327548
      WHEN 1709 => Ti := "000001010100010101110010111110101001101111100110"; --    +345458    -353306
      WHEN 1710 => Ti := "111110101011011011001001111001110011110000010101"; --    -346423   -1623019
      WHEN 1711 => Ti := "000010000101100101000111111101101110111001000101"; --    +547143    -594363
      WHEN 1712 => Ti := "000011000001011001001100111110001001010110111110"; --    +792140    -485954
      WHEN 1713 => Ti := "111111100101110010101011000010100011101000010000"; --    -107349    +670224
      WHEN 1714 => Ti := "111010111110011100111111000000101101010111011111"; --   -1317057    +185823
      WHEN 1715 => Ti := "000101010000001001000111000000100110010100000101"; --   +1376839    +156933
      WHEN 1716 => Ti := "111101001010101001110111111101110100010000111111"; --    -742793    -572353
      WHEN 1717 => Ti := "111011001011000100000101111110011000010011001010"; --   -1265403    -424758
      WHEN 1718 => Ti := "111111110110000101101010000000110000001001011101"; --     -40598    +197213
      WHEN 1719 => Ti := "001000101111110001000101111101111101011101111000"; --   +2292805    -534664
      WHEN 1720 => Ti := "000010001000001000101011000000001101000111110111"; --    +557611     +53751
      WHEN 1721 => Ti := "000010000000010101000101111101010100110111100010"; --    +525637    -700958
      WHEN 1722 => Ti := "111111011110000001010001111110010101111000100010"; --    -139183    -434654
      WHEN 1723 => Ti := "000000100000000100000001111001100100011111011010"; --    +131329   -1685542
      WHEN 1724 => Ti := "111100110111011010010001111101101011001101100110"; --    -821615    -609434
      WHEN 1725 => Ti := "000011100111000000110001000000110101011000111100"; --    +946225    +218684
      WHEN 1726 => Ti := "000000010101010001101101000001011111000001101101"; --     +87149    +389229
      WHEN 1727 => Ti := "111101010111100000101100111110001100000100010110"; --    -690132    -474858
      WHEN 1728 => Ti := "000001110010011110100010000011010101101000011001"; --    +468898    +875033
      WHEN 1729 => Ti := "111011111011000000101110111111111001111101101011"; --   -1069010     -24725
      WHEN 1730 => Ti := "000011000100100000100111111110110001010001001100"; --    +804903    -322484
      WHEN 1731 => Ti := "000001001101100001101000111111001001001000110110"; --    +317544    -224714
      WHEN 1732 => Ti := "000001100110010000010111111111101001011100001100"; --    +418839     -92404
      WHEN 1733 => Ti := "000101000111111010001110000010001100111010110001"; --   +1343118    +577201
      WHEN 1734 => Ti := "000000011001000110010010111101110001011111110101"; --    +102802    -583691
      WHEN 1735 => Ti := "111111010110110111010010111110101101111101101111"; --    -168494    -336017
      WHEN 1736 => Ti := "111110101011101010100001111101111010110100011001"; --    -345439    -545511
      WHEN 1737 => Ti := "111100111011011110010000111111000100100111110010"; --    -804976    -243214
      WHEN 1738 => Ti := "000001110111010011100101000000010101001100101000"; --    +488677     +86824
      WHEN 1739 => Ti := "000001011011101101001000000001100100000100011011"; --    +375624    +409883
      WHEN 1740 => Ti := "111110000110111101100110111111001111000101110011"; --    -495770    -200333
      WHEN 1741 => Ti := "000100100100100110001011111011011001000010011101"; --   +1198475   -1208163
      WHEN 1742 => Ti := "111001101101001011111001111111010111010111101000"; --   -1649927    -166424
      WHEN 1743 => Ti := "000000111001101010111111000001001010000110101010"; --    +236223    +303530
      WHEN 1744 => Ti := "111110101001011101100100111111110000100001011000"; --    -354460     -63400
      WHEN 1745 => Ti := "000000111000111100111111111110110000011011010100"; --    +233279    -325932
      WHEN 1746 => Ti := "000011011000000001110111111110111000001010010100"; --    +884855    -294252
      WHEN 1747 => Ti := "000010110100110111010000111111110101111100001010"; --    +740816     -41206
      WHEN 1748 => Ti := "111110101001110010111110000111010011110000111110"; --    -353090   +1915966
      WHEN 1749 => Ti := "111101110010101001000001111111111001111111111000"; --    -579007     -24584
      WHEN 1750 => Ti := "111100001001101001011000000000010001001001100110"; --   -1009064     +70246
      WHEN 1751 => Ti := "111101010101000010110011000000001101101000100100"; --    -700237     +55844
      WHEN 1752 => Ti := "000010001100100100101000111101011011110000100100"; --    +575784    -672732
      WHEN 1753 => Ti := "111111100000010001100000000011010001100101111110"; --    -129952    +858494
      WHEN 1754 => Ti := "111110100111000001011011000000001001000110101111"; --    -364453     +37295
      WHEN 1755 => Ti := "111100011011001101110101111100001101001111000010"; --    -937099    -994366
      WHEN 1756 => Ti := "111111000011011100011110000000000011111100111110"; --    -248034     +16190
      WHEN 1757 => Ti := "000000111110111011010111000011101110111101011011"; --    +257751    +978779
      WHEN 1758 => Ti := "000001111100010000111001000000011011101010011101"; --    +508985    +113309
      WHEN 1759 => Ti := "111010110101010111110100000000010011010111111110"; --   -1354252     +79358
      WHEN 1760 => Ti := "000000001010011010110010111100000000001110010010"; --     +42674   -1047662
      WHEN 1761 => Ti := "111111101001011001011001000000001011110011011000"; --     -92583     +48344
      WHEN 1762 => Ti := "111100111110010101101110000010000101000010110011"; --    -793234    +544947
      WHEN 1763 => Ti := "111111101100001011101011111011100010110101101000"; --     -81173   -1168024
      WHEN 1764 => Ti := "000000100101010001011000111110000100111111000111"; --    +152664    -503865
      WHEN 1765 => Ti := "000001111111000010000001111110101111110010101111"; --    +520321    -328529
      WHEN 1766 => Ti := "000001111110011111000100000011011110011101100010"; --    +518084    +911202
      WHEN 1767 => Ti := "111110111101101000101010111111011100110100000010"; --    -271830    -144126
      WHEN 1768 => Ti := "111110100111101011010101000100010001110100000001"; --    -361771   +1121537
      WHEN 1769 => Ti := "111111110011111111101111000011110000001010100010"; --     -49169    +983714
      WHEN 1770 => Ti := "111011011101100010110100111110110100011101000110"; --   -1189708    -309434
      WHEN 1771 => Ti := "111101110000010011100101111011010101100010011111"; --    -588571   -1222497
      WHEN 1772 => Ti := "000000001100000000110010000001010111100010111010"; --     +49202    +358586
      WHEN 1773 => Ti := "000100001010110100010011111110100000111110100101"; --   +1092883    -389211
      WHEN 1774 => Ti := "111111001001111111110000111100011101000101111110"; --    -221200    -929410
      WHEN 1775 => Ti := "111011100110101110101111111101000001111011000111"; --   -1152081    -778553
      WHEN 1776 => Ti := "000010000100100010010001000000110011010100111111"; --    +542865    +210239
      WHEN 1777 => Ti := "111010111001100101101001111110111010111100010011"; --   -1336983    -282861
      WHEN 1778 => Ti := "000001101011001000111001111111001010111100000001"; --    +438841    -217343
      WHEN 1779 => Ti := "111110010001101110000111000000001001010011111111"; --    -451705     +38143
      WHEN 1780 => Ti := "111110011101011101010101000001000101001111100010"; --    -403627    +283618
      WHEN 1781 => Ti := "000010101001001001100011000001010010010101010001"; --    +692835    +337233
      WHEN 1782 => Ti := "000001011010111010111001111100101000100100001000"; --    +372409    -882424
      WHEN 1783 => Ti := "000010000110110000000101111101100110110001100110"; --    +551941    -627610
      WHEN 1784 => Ti := "111100001111100010000111111110000001111011110110"; --    -984953    -516362
      WHEN 1785 => Ti := "111110110110101100101010111110110000110001001111"; --    -300246    -324529
      WHEN 1786 => Ti := "111111101111010100011011111100000110110001000101"; --     -68325   -1020859
      WHEN 1787 => Ti := "111011100000111101101111000010110110001010110111"; --   -1175697    +746167
      WHEN 1788 => Ti := "000010011000000101111100111101010010011000101110"; --    +622972    -711122
      WHEN 1789 => Ti := "111111110010101111000000000000011011101100111010"; --     -54336    +113466
      WHEN 1790 => Ti := "111011111110001100100001000000000010101101101011"; --   -1055967     +11115
      WHEN 1791 => Ti := "111101010111001010110010111101110010100111110001"; --    -691534    -579087
      WHEN 1792 => Ti := "000100100111111101001000000100001110001010010101"; --   +1212232   +1106581
      WHEN 1793 => Ti := "000000001001111110000011111111010000001010111110"; --     +40835    -195906
      WHEN 1794 => Ti := "000001110100011100111111111101100111011011101111"; --    +476991    -624913
      WHEN 1795 => Ti := "111100111110001010011101111011110111010101011001"; --    -793955   -1084071
      WHEN 1796 => Ti := "111100111111110100010000111110100010001100101000"; --    -787184    -384216
      WHEN 1797 => Ti := "111100110011101000101000111111110010001111000100"; --    -837080     -56380
      WHEN 1798 => Ti := "000011000100101100100110111111001011100011000011"; --    +805670    -214845
      WHEN 1799 => Ti := "111011110011100001110101111111000100111110100100"; --   -1099659    -241756
      WHEN 1800 => Ti := "111011011100100100101100111101001100011111101101"; --   -1193684    -735251
      WHEN 1801 => Ti := "111111111001001100100111111101001110011101100101"; --     -27865    -727195
      WHEN 1802 => Ti := "111111111010010010101110000010000010001100010001"; --     -23378    +533265
      WHEN 1803 => Ti := "000011111100001101110001111010101000100010101011"; --   +1033073   -1406805
      WHEN 1804 => Ti := "111011111000100111000100000000000100110000000010"; --   -1078844     +19458
      WHEN 1805 => Ti := "000001010001110000011011000010001100001011001001"; --    +334875    +574153
      WHEN 1806 => Ti := "111011011000101111101100111011110100001001001101"; --   -1209364   -1097139
      WHEN 1807 => Ti := "111110101101110000000001111101010101010101000100"; --    -336895    -699068
      WHEN 1808 => Ti := "000000111101000010010110000011001110110111010011"; --    +250006    +847315
      WHEN 1809 => Ti := "000000000010101010111001000000101010011111011011"; --     +10937    +174043
      WHEN 1810 => Ti := "000010100011010000010001111101111000101100100101"; --    +668689    -554203
      WHEN 1811 => Ti := "000001000000101100100011000000010110111100100100"; --    +264995     +93988
      WHEN 1812 => Ti := "000001111110101000111011111110111100011111111100"; --    +518715    -276484
      WHEN 1813 => Ti := "000001001000100100101010111110001101111110010001"; --    +297258    -467055
      WHEN 1814 => Ti := "000000101100111001111101111110101000100111101010"; --    +183933    -357910
      WHEN 1815 => Ti := "000100101011010010001000000110001101101000111100"; --   +1225864   +1628732
      WHEN 1816 => Ti := "000001010101111010011011111111001100010010100010"; --    +351899    -211806
      WHEN 1817 => Ti := "000000001000111000100101000001001001111010011001"; --     +36389    +302745
      WHEN 1818 => Ti := "111110001011111100101100000010111111001000110111"; --    -475348    +782903
      WHEN 1819 => Ti := "111101111000000000011000111010101010110001100110"; --    -557032   -1397658
      WHEN 1820 => Ti := "111111010110100011011011111100011100000010010100"; --    -169765    -933740
      WHEN 1821 => Ti := "111110001011001011011011111110010001110101110011"; --    -478501    -451213
      WHEN 1822 => Ti := "000011000111110111001001000011001110011000110111"; --    +818633    +845367
      WHEN 1823 => Ti := "111110010100101001110011000000010101100101010011"; --    -439693     +88403
      WHEN 1824 => Ti := "111011000101011011010100000011000011100111010011"; --   -1288492    +801235
      WHEN 1825 => Ti := "111110000101101110001101000001100011111100000100"; --    -500851    +409348
      WHEN 1826 => Ti := "111101010011011101100100000010100100101011011101"; --    -706716    +674525
      WHEN 1827 => Ti := "111110111100001001001100000010000010001110010110"; --    -277940    +533398
      WHEN 1828 => Ti := "000000011011001101011110000011101010111101010000"; --    +111454    +962384
      WHEN 1829 => Ti := "000010111111001001010101111111010011111100011000"; --    +782933    -180456
      WHEN 1830 => Ti := "111010101100000010110111111110100011101110000101"; --   -1392457    -377979
      WHEN 1831 => Ti := "111100010001111100011111111011101000010110011101"; --    -975073   -1145443
      WHEN 1832 => Ti := "000000111011100000000011000001011100001000001000"; --    +243715    +377352
      WHEN 1833 => Ti := "000000101100111001100101111110011100111100000001"; --    +183909    -405759
      WHEN 1834 => Ti := "111111000110111001110110000001010110100001010101"; --    -233866    +354389
      WHEN 1835 => Ti := "000001000111110010000010000010100000110110011011"; --    +294018    +658843
      WHEN 1836 => Ti := "000100100001010000111011111110110000101000000001"; --   +1184827    -325119
      WHEN 1837 => Ti := "000001011110111011011100000001001100000101110011"; --    +388828    +311667
      WHEN 1838 => Ti := "000000111111111001101100111101000100100000011010"; --    +261740    -767974
      WHEN 1839 => Ti := "111100111101100001000111000010110011000101010001"; --    -796601    +733521
      WHEN 1840 => Ti := "000011101001110010011100111110000101001101000000"; --    +957596    -502976
      WHEN 1841 => Ti := "111000101011101010011000111100011101011111101110"; --   -1918312    -927762
      WHEN 1842 => Ti := "111101011101011010010110000100111010101010001001"; --    -665962   +1288841
      WHEN 1843 => Ti := "111111010011011000000011111110100111001011111010"; --    -182781    -363782
      WHEN 1844 => Ti := "111101011110110000010101000000111001111001010111"; --    -660459    +237143
      WHEN 1845 => Ti := "111111110001001100001110000011000110101001000010"; --     -60658    +813634
      WHEN 1846 => Ti := "111100100011011001001010111111100001110010101010"; --    -903606    -123734
      WHEN 1847 => Ti := "000001000110110111110000111011111010111011110111"; --    +290288   -1069321
      WHEN 1848 => Ti := "111101111100100100111100000000101111111111000010"; --    -538308    +196546
      WHEN 1849 => Ti := "111101000001110110100010000000110111110000001110"; --    -778846    +228366
      WHEN 1850 => Ti := "111100111000100000110111111110110000000101111001"; --    -817097    -327303
      WHEN 1851 => Ti := "000001110000100001011101000000101100111110100001"; --    +460893    +184225
      WHEN 1852 => Ti := "000011101010010100000000000001111011101010110111"; --    +959744    +506551
      WHEN 1853 => Ti := "111101110101110101001111111111011110011011011111"; --    -565937    -137505
      WHEN 1854 => Ti := "000011011110000110010010111011100101001101100100"; --    +909714   -1158300
      WHEN 1855 => Ti := "000010110010001111010110111101000100101101111001"; --    +730070    -767111
      WHEN 1856 => Ti := "111010110010110100111111111101001000110011100100"; --   -1364673    -750364
      WHEN 1857 => Ti := "111110010000100010000101111111100111011101110010"; --    -456571    -100494
      WHEN 1858 => Ti := "111110001001001110101100111100110100100001111101"; --    -486484    -833411
      WHEN 1859 => Ti := "000010010100101000101010111101010000011100001011"; --    +608810    -719093
      WHEN 1860 => Ti := "000000001110101110101110000010011101111010101100"; --     +60334    +646828
      WHEN 1861 => Ti := "000010000110110100110000000000011111001010101100"; --    +552240    +127660
      WHEN 1862 => Ti := "111110010100011111101000000011001001101000001011"; --    -440344    +825867
      WHEN 1863 => Ti := "000000000010011010010011111101110100011001001110"; --      +9875    -571826
      WHEN 1864 => Ti := "000001000010010110101100111100010101001101000101"; --    +271788    -961723
      WHEN 1865 => Ti := "111111001001000110001011000011110010010101011000"; --    -224885    +992600
      WHEN 1866 => Ti := "111101110111110011111000111101111000010000110101"; --    -557832    -555979
      WHEN 1867 => Ti := "111111010111001001100111111111001001000011111011"; --    -167321    -225029
      WHEN 1868 => Ti := "111001111110111111010001111110010110010110111000"; --   -1577007    -432712
      WHEN 1869 => Ti := "000001011010010001100011000000010010101001111011"; --    +369763     +76411
      WHEN 1870 => Ti := "000000110000001010111100000001100110111111011011"; --    +197308    +421851
      WHEN 1871 => Ti := "111101101111110101001011111111000100101000101010"; --    -590517    -243158
      WHEN 1872 => Ti := "000010011010100111100000000000101010101110010110"; --    +633312    +174998
      WHEN 1873 => Ti := "000011101110101110100110000100010011001000011111"; --    +977830   +1126943
      WHEN 1874 => Ti := "000001011001011010000000000001000111101101100101"; --    +366208    +293733
      WHEN 1875 => Ti := "000001011010001100010011000000110001110001100111"; --    +369427    +203879
      WHEN 1876 => Ti := "111110110111001100110000000000010010001101101111"; --    -298192     +74607
      WHEN 1877 => Ti := "111110111010101100111011111101110100111100001001"; --    -283845    -569591
      WHEN 1878 => Ti := "000001011100001010111101111011111111010001001101"; --    +377533   -1051571
      WHEN 1879 => Ti := "000000000111100111100000000010001110001010100011"; --     +31200    +582307
      WHEN 1880 => Ti := "000000011111000101010111111101010011100011011101"; --    +127319    -706339
      WHEN 1881 => Ti := "000011000000010101011001111101111010001000101001"; --    +787801    -548311
      WHEN 1882 => Ti := "111111110001000011001011111111110100110100110101"; --     -61237     -45771
      WHEN 1883 => Ti := "111001111010011100010110000011000111000100110010"; --   -1595626    +815410
      WHEN 1884 => Ti := "000001101111000011110101111110111100011111111101"; --    +454901    -276483
      WHEN 1885 => Ti := "000010010001000101111100000001010011110001111101"; --    +594300    +343165
      WHEN 1886 => Ti := "000010010101100000110011111100000010101110101100"; --    +612403   -1037396
      WHEN 1887 => Ti := "000011100011011001011010000011000110100101010011"; --    +931418    +813395
      WHEN 1888 => Ti := "111100101100110111010110111111010101011000011000"; --    -864810    -174568
      WHEN 1889 => Ti := "111110101010011111110100000001010101000001000110"; --    -350220    +348230
      WHEN 1890 => Ti := "111111010000101101100001111011011010101100010011"; --    -193695   -1201389
      WHEN 1891 => Ti := "000000111001110111110100111111011101010111111000"; --    +237044    -141832
      WHEN 1892 => Ti := "000000110100101101100000000010111000011101000111"; --    +215904    +755527
      WHEN 1893 => Ti := "111111100111000000000111000101111011000110101100"; --    -102393   +1552812
      WHEN 1894 => Ti := "000001000011001110000110111101000110000010000110"; --    +275334    -761722
      WHEN 1895 => Ti := "000001101100010011000100000001110000011001011010"; --    +443588    +460378
      WHEN 1896 => Ti := "000010101011101101111011111100000101011111101010"; --    +703355   -1026070
      WHEN 1897 => Ti := "111110010101000000110110000001011011101101100010"; --    -438218    +375650
      WHEN 1898 => Ti := "111111001010011110011110111111001010011101010001"; --    -219234    -219311
      WHEN 1899 => Ti := "000010111001110111110111000010101100011100100001"; --    +761335    +706337
      WHEN 1900 => Ti := "111111101111101000110101111101010111100101111111"; --     -67019    -689793
      WHEN 1901 => Ti := "111111011011111101101111111010100100100010000011"; --    -147601   -1423229
      WHEN 1902 => Ti := "111111011011001001000000111111110001010010011100"; --    -150976     -60260
      WHEN 1903 => Ti := "111011000010101110110101111101011000000010001111"; --   -1299531    -687985
      WHEN 1904 => Ti := "000011001011000101011001111010111101000101110101"; --    +831833   -1322635
      WHEN 1905 => Ti := "000000001010010101010110000001001010100101100101"; --     +42326    +305509
      WHEN 1906 => Ti := "111100010111100001111101000011000110001111110100"; --    -952195    +812020
      WHEN 1907 => Ti := "111101111001001110100011111011001111000000001101"; --    -552029   -1249267
      WHEN 1908 => Ti := "000000101111011000101010111101011110111011101101"; --    +194090    -659731
      WHEN 1909 => Ti := "111101011011101001110110111100011010000100110011"; --    -673162    -941773
      WHEN 1910 => Ti := "111100101001101011111101111110010100110001011000"; --    -877827    -439208
      WHEN 1911 => Ti := "111111001100001011101100000001001110000001001110"; --    -212244    +319566
      WHEN 1912 => Ti := "000100110100111110100110111100111111100111111110"; --   +1265574    -787970
      WHEN 1913 => Ti := "000000001000101011100100000000001101000001110000"; --     +35556     +53360
      WHEN 1914 => Ti := "111100111001000001111000000001100100101111100011"; --    -814984    +412643
      WHEN 1915 => Ti := "000001000011100001010111000000110100011010110111"; --    +276567    +214711
      WHEN 1916 => Ti := "000010100011111101001000000000011110011010111101"; --    +671560    +124605
      WHEN 1917 => Ti := "111110011010110010101010111110010011100110111000"; --    -414550    -443976
      WHEN 1918 => Ti := "000100001100010010100011111011111101000010100000"; --   +1098915   -1060704
      WHEN 1919 => Ti := "111111000101100000011010000001001110101100011001"; --    -239590    +322329
      WHEN 1920 => Ti := "111101001111110011110110000001011100111001010101"; --    -721674    +380501
      WHEN 1921 => Ti := "000011110000010001011111111101001011000011111100"; --    +984159    -741124
      WHEN 1922 => Ti := "000011111001101001111110111111100011111101011110"; --   +1022590    -114850
      WHEN 1923 => Ti := "000001001011011100011010111101001001101001101100"; --    +309018    -746900
      WHEN 1924 => Ti := "111111000010000100111000111110000111110101000011"; --    -253640    -492221
      WHEN 1925 => Ti := "111111111000111101110000111100011010101011000010"; --     -28816    -939326
      WHEN 1926 => Ti := "111010001101100100010111111110011101011001111101"; --   -1517289    -403843
      WHEN 1927 => Ti := "000011101011111010011000111111011100010110100010"; --    +966296    -146014
      WHEN 1928 => Ti := "000011010001010000100100000001010000110000010101"; --    +857124    +330773
      WHEN 1929 => Ti := "111111010010100011010001000010010001011011000000"; --    -186159    +595648
      WHEN 1930 => Ti := "000001101100100000100101111010101000001111001111"; --    +444453   -1408049
      WHEN 1931 => Ti := "111101011011001001110011111101010100000110000000"; --    -675213    -704128
      WHEN 1932 => Ti := "000001101001001111111101000011001110110101110110"; --    +431101    +847222
      WHEN 1933 => Ti := "000010111110011000100111111110001010101001011110"; --    +779815    -480674
      WHEN 1934 => Ti := "111111111000010001011101111110110111000111101111"; --     -31651    -298513
      WHEN 1935 => Ti := "000101100101010010111000000000001100110101000110"; --   +1463480     +52550
      WHEN 1936 => Ti := "000010101100001010010100000001110010001000110111"; --    +705172    +467511
      WHEN 1937 => Ti := "111100010010010011110111000001111111110010110010"; --    -973577    +523442
      WHEN 1938 => Ti := "111111010100000000011111111101111001110001101010"; --    -180193    -549782
      WHEN 1939 => Ti := "111101101110001100101001000000110100001011101111"; --    -597207    +213743
      WHEN 1940 => Ti := "000000000101101001111010000000001000100101001000"; --     +23162     +35144
      WHEN 1941 => Ti := "000011100000001100100111000100100111110011111000"; --    +918311   +1211640
      WHEN 1942 => Ti := "000001011110010101110100111111010110100000111111"; --    +386420    -169921
      WHEN 1943 => Ti := "111101001101101111001100111110110100000010101111"; --    -730164    -311121
      WHEN 1944 => Ti := "000010011111011011110010111110111000010111000000"; --    +653042    -293440
      WHEN 1945 => Ti := "111111000010110000011010000011100001100001000111"; --    -250854    +923719
      WHEN 1946 => Ti := "000100011110101110000010111111011111110010000101"; --   +1174402    -131963
      WHEN 1947 => Ti := "111100100110110100010011000000101011000000100000"; --    -889581    +176160
      WHEN 1948 => Ti := "000000100011100100001001111101110011111100101010"; --    +145673    -573654
      WHEN 1949 => Ti := "111110001001100110101011000000111110011101000010"; --    -484949    +255810
      WHEN 1950 => Ti := "000001101010001001101110111111011110000011111111"; --    +434798    -139009
      WHEN 1951 => Ti := "000011011001000000111100000011100110110111010011"; --    +888892    +945619
      WHEN 1952 => Ti := "000010110101011010011010000010010100110000100011"; --    +743066    +609315
      WHEN 1953 => Ti := "000010101101100110001110000010110000111000100001"; --    +711054    +724513
      WHEN 1954 => Ti := "111110000011100111001110111011110111000111111010"; --    -509490   -1084934
      WHEN 1955 => Ti := "000000110110110100011010000010001110000011111001"; --    +224538    +581881
      WHEN 1956 => Ti := "111100001100010111111001111110100001000111001010"; --    -997895    -388662
      WHEN 1957 => Ti := "111111000110000101000011000001000111000100001011"; --    -237245    +291083
      WHEN 1958 => Ti := "111110010010011011000011000001011111110110110110"; --    -448829    +392630
      WHEN 1959 => Ti := "000000111100011111011001000000100011000101000001"; --    +247769    +143681
      WHEN 1960 => Ti := "000011011111100010101110000011101000001011111101"; --    +915630    +951037
      WHEN 1961 => Ti := "000000111100010000110111000001010100010001111101"; --    +246839    +345213
      WHEN 1962 => Ti := "000001011001101111001010000010110100010110011000"; --    +367562    +738712
      WHEN 1963 => Ti := "111011000010101010001101000001110111111000110011"; --   -1299827    +491059
      WHEN 1964 => Ti := "000000000100111001000100111101010011000100001010"; --     +20036    -708342
      WHEN 1965 => Ti := "000000100111000010010011111110110101110001101111"; --    +159891    -304017
      WHEN 1966 => Ti := "000001001101000101111101000010000010101000000100"; --    +315773    +535044
      WHEN 1967 => Ti := "000100001110011001100000000010111111010110011011"; --   +1107552    +783771
      WHEN 1968 => Ti := "000000101010101110011010000001101011000100000100"; --    +175002    +438532
      WHEN 1969 => Ti := "111111001100111000110010111101011100000010000010"; --    -209358    -671614
      WHEN 1970 => Ti := "111011100101000101101011000010010110010001110100"; --   -1158805    +615540
      WHEN 1971 => Ti := "000000101110111001001100000010101010011011111110"; --    +192076    +698110
      WHEN 1972 => Ti := "111110000110011011100101111101111011000001001101"; --    -497947    -544691
      WHEN 1973 => Ti := "000111010101111010111101111110100111010011101111"; --   +1924797    -363281
      WHEN 1974 => Ti := "111101101010001001001100111101111000000111011100"; --    -613812    -556580
      WHEN 1975 => Ti := "111111110111010010000111000001010000110100010101"; --     -35705    +331029
      WHEN 1976 => Ti := "000011000010001011010101111110011111001100101101"; --    +795349    -396499
      WHEN 1977 => Ti := "111111000101000100110001000000110010010000001011"; --    -241359    +205835
      WHEN 1978 => Ti := "111100110011000100100110000010111110111110000110"; --    -839386    +782214
      WHEN 1979 => Ti := "111100101111111011010100111101110110000110001101"; --    -852268    -564851
      WHEN 1980 => Ti := "000010001000010100110101000011010010111110111001"; --    +558389    +864185
      WHEN 1981 => Ti := "111110001100011100100111111111000101010001011111"; --    -473305    -240545
      WHEN 1982 => Ti := "111100110101001110001001111111111101100011011101"; --    -830583     -10019
      WHEN 1983 => Ti := "000100111000111000001101000001000000111010111001"; --   +1281549    +265913
      WHEN 1984 => Ti := "000000111010001100110101000110111100111011000011"; --    +238389   +1822403
      WHEN 1985 => Ti := "111011001101111001010000000010101111110010101001"; --   -1253808    +720041
      WHEN 1986 => Ti := "111110010110010101001111111100011010111101000011"; --    -432817    -938173
      WHEN 1987 => Ti := "111111001111011111110000111100110111001101110011"; --    -198672    -822413
      WHEN 1988 => Ti := "111110001010110001010100000010110001001110110100"; --    -480172    +725940
      WHEN 1989 => Ti := "000011111010000100100100000010101100001010011001"; --   +1024292    +705177
      WHEN 1990 => Ti := "111111110110001110101101111010011000010000011101"; --     -40019   -1473507
      WHEN 1991 => Ti := "111101001111010010100111111110111100101011101001"; --    -723801    -275735
      WHEN 1992 => Ti := "111101011100000100001000111111110111111000100101"; --    -671480     -33243
      WHEN 1993 => Ti := "000100110001110011010001000000100111111000010010"; --   +1252561    +163346
      WHEN 1994 => Ti := "000001100101101110100101000000100000000010100001"; --    +416677    +131233
      WHEN 1995 => Ti := "111101101111110110110101000001010111111100011010"; --    -590411    +360218
      WHEN 1996 => Ti := "111110111010101100011110111111100101111110000000"; --    -283874    -106624
      WHEN 1997 => Ti := "000001011001000111011100111100101010010111000010"; --    +365020    -875070
      WHEN 1998 => Ti := "111101011000001101110110000001100011000100100100"; --    -687242    +405796
      WHEN 1999 => Ti := "000010000001100011011101111110100101000011100000"; --    +530653    -372512
      WHEN 2000 => Ti := "111011110101111101011101111110000110001110011010"; --   -1089699    -498790
      WHEN 2001 => Ti := "111100010001011001101101000011011000110110111001"; --    -977299    +888249
      WHEN 2002 => Ti := "000000010100001101011000111110100111000001011011"; --     +82776    -364453
      WHEN 2003 => Ti := "000001010011010000101011111101100011100100110011"; --    +341035    -640717
      WHEN 2004 => Ti := "000001001100001010010010000001000110000011101101"; --    +311954    +286957
      WHEN 2005 => Ti := "000001000000101101111000000010100101000001010111"; --    +265080    +675927
      WHEN 2006 => Ti := "111111010110111110101010111011101001100101101100"; --    -168022   -1140372
      WHEN 2007 => Ti := "000000100000011101011111111110000000101100010011"; --    +132959    -521453
      WHEN 2008 => Ti := "000000000100010101111111111110010011000010100000"; --     +17791    -446304
      WHEN 2009 => Ti := "000010111100100110100101111010000000101101000010"; --    +772517   -1569982
      WHEN 2010 => Ti := "000000100100101110100000000100111000001011100011"; --    +150432   +1278691
      WHEN 2011 => Ti := "111110100100101000001101111100000011111000001010"; --    -374259   -1032694
      WHEN 2012 => Ti := "000010000001100100010111000000001000110111101100"; --    +530711     +36332
      WHEN 2013 => Ti := "000001110010011000011111111101110110100010101111"; --    +468511    -563025
      WHEN 2014 => Ti := "111110010010100100000001000000101100111011001010"; --    -448255    +184010
      WHEN 2015 => Ti := "111111101011010011111001000000011101010001100110"; --     -84743    +119910
      WHEN 2016 => Ti := "000010001100111011101101111111011100111010100100"; --    +577261    -143708
      WHEN 2017 => Ti := "000001010001001000111101000000100100001001000010"; --    +332349    +148034
      WHEN 2018 => Ti := "111110011001001111111011000011111010010100110001"; --    -420869   +1025329
      WHEN 2019 => Ti := "000001010010101110101001000000110111010100001111"; --    +338857    +226575
      WHEN 2020 => Ti := "111110111100000101101100111111010011001100010010"; --    -278164    -183534
      WHEN 2021 => Ti := "111011001110011111100010111010101000100000011100"; --   -1251358   -1406948
      WHEN 2022 => Ti := "000011001101100101111000111111000101011010011001"; --    +842104    -239975
      WHEN 2023 => Ti := "000001001011101011111110000010100000111111101011"; --    +310014    +659435
      WHEN 2024 => Ti := "111100101011101100110101111110110110011000100000"; --    -869579    -301536
      WHEN 2025 => Ti := "111111011101010011101001000010011100100110110001"; --    -142103    +641457
      WHEN 2026 => Ti := "111111000110110101111110111101001101100100011001"; --    -234114    -730855
      WHEN 2027 => Ti := "111011000010011010111010111110101111010111010100"; --   -1300806    -330284
      WHEN 2028 => Ti := "000100001010111101000011111111011110100111101011"; --   +1093443    -136725
      WHEN 2029 => Ti := "000000001000000001111011000011000010000110001010"; --     +32891    +795018
      WHEN 2030 => Ti := "000001101010001110011001000001001010110011001010"; --    +435097    +306378
      WHEN 2031 => Ti := "111111000001110010110011111100100001111010101000"; --    -254797    -909656
      WHEN 2032 => Ti := "000001001101101111101100000001011011110000110110"; --    +318444    +375862
      WHEN 2033 => Ti := "000011010110111001100000000001001101000111110111"; --    +880224    +315895
      WHEN 2034 => Ti := "000010011101100000101101000000110100110110000010"; --    +645165    +216450
      WHEN 2035 => Ti := "000000101011100011100011111110011010011000000010"; --    +178403    -416254
      WHEN 2036 => Ti := "111111000111111100000101111100100101000100000000"; --    -229627    -896768
      WHEN 2037 => Ti := "111110100000000000011001111100111000101100111110"; --    -393191    -816322
      WHEN 2038 => Ti := "111111110001111000000100000110100100001010001011"; --     -57852   +1720971
      WHEN 2039 => Ti := "000001101000111110100010111111001101111001011110"; --    +429986    -205218
      WHEN 2040 => Ti := "000000101111011100010001111111000011101111100000"; --    +194321    -246816
      WHEN 2041 => Ti := "000011101010010111011101111111010000010010101010"; --    +959965    -195414
      WHEN 2042 => Ti := "000000000100000000111000111101101010101101110011"; --     +16440    -611469
      WHEN 2043 => Ti := "111101101101001010011111000010101000000000011100"; --    -601441    +688156
      WHEN 2044 => Ti := "111110111001011010100111000101110001110110111101"; --    -289113   +1514941
      WHEN 2045 => Ti := "111011011111101001010110111111001110000111101011"; --   -1181098    -204309
      WHEN 2046 => Ti := "000000010011010111110000111110101101110010011010"; --     +79344    -336742
      WHEN 2047 => Ti := "000010111100110010111101000000001100010100111001"; --    +773309     +50489
      WHEN OTHERS => NULL;
    END CASE; 
    T <= Ti; 
  END PROCESS; 
END ARCHITECTURE arch_rom; 



