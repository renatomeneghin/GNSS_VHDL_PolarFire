-- CoreDDS Output Golden Test Vectors.
-- Test run length = 510

LIBRARY IEEE; 
  USE IEEE.std_logic_1164.all; 

ENTITY dds_bhvTestVectOut IS
  GENERIC ( OUTPUT_BITS    : INTEGER := 10  );
  PORT  ( sample_num       :  IN integer;
          goldSin, goldCos : OUT STD_LOGIC_VECTOR(OUTPUT_BITS-1 DOWNTO 0) );
END ENTITY dds_bhvTestVectOut;

ARCHITECTURE rtl of dds_bhvTestVectOut IS
  BEGIN
    PROCESS (sample_num)
      BEGIN
        CASE sample_num IS
          WHEN   0 => goldSin <= "111111111111";
                      goldCos <= "010000000000";
          WHEN   1 => goldSin <= "111111111111";
                      goldCos <= "010000000000";
          WHEN   2 => goldSin <= "111110011011";
                      goldCos <= "001111111011";
          WHEN   3 => goldSin <= "111100110111";
                      goldCos <= "001111101100";
          WHEN   4 => goldSin <= "111011010110";
                      goldCos <= "001111010100";
          WHEN   5 => goldSin <= "111001110111";
                      goldCos <= "001110110010";
          WHEN   6 => goldSin <= "111000011101";
                      goldCos <= "001110000111";
          WHEN   7 => goldSin <= "110111000110";
                      goldCos <= "001101010011";
          WHEN   8 => goldSin <= "110101110110";
                      goldCos <= "001100010111";
          WHEN   9 => goldSin <= "110100101011";
                      goldCos <= "001011010100";
          WHEN  10 => goldSin <= "110011101000";
                      goldCos <= "001010001001";
          WHEN  11 => goldSin <= "110010101100";
                      goldCos <= "001000111000";
          WHEN  12 => goldSin <= "110001111001";
                      goldCos <= "000111100010";
          WHEN  13 => goldSin <= "110001001110";
                      goldCos <= "000110000111";
          WHEN  14 => goldSin <= "110000101100";
                      goldCos <= "000100101000";
          WHEN  15 => goldSin <= "110000010100";
                      goldCos <= "000011000111";
          WHEN  16 => goldSin <= "110000000101";
                      goldCos <= "000001100100";
          WHEN  17 => goldSin <= "110000000000";
                      goldCos <= "111111111111";
          WHEN  18 => goldSin <= "110000000101";
                      goldCos <= "111110011011";
          WHEN  19 => goldSin <= "110000010100";
                      goldCos <= "111100110111";
          WHEN  20 => goldSin <= "110000101100";
                      goldCos <= "111011010110";
          WHEN  21 => goldSin <= "110001001110";
                      goldCos <= "111001110111";
          WHEN  22 => goldSin <= "110001111001";
                      goldCos <= "111000011101";
          WHEN  23 => goldSin <= "110010101101";
                      goldCos <= "110111000110";
          WHEN  24 => goldSin <= "110011101001";
                      goldCos <= "110101110110";
          WHEN  25 => goldSin <= "110100101100";
                      goldCos <= "110100101011";
          WHEN  26 => goldSin <= "110101110111";
                      goldCos <= "110011101000";
          WHEN  27 => goldSin <= "110111001000";
                      goldCos <= "110010101100";
          WHEN  28 => goldSin <= "111000011110";
                      goldCos <= "110001111001";
          WHEN  29 => goldSin <= "111001111001";
                      goldCos <= "110001001110";
          WHEN  30 => goldSin <= "111011011000";
                      goldCos <= "110000101100";
          WHEN  31 => goldSin <= "111100111001";
                      goldCos <= "110000010100";
          WHEN  32 => goldSin <= "111110011100";
                      goldCos <= "110000000101";
          WHEN  33 => goldSin <= "000000000001";
                      goldCos <= "110000000000";
          WHEN  34 => goldSin <= "000001100101";
                      goldCos <= "110000000101";
          WHEN  35 => goldSin <= "000011001001";
                      goldCos <= "110000010100";
          WHEN  36 => goldSin <= "000100101010";
                      goldCos <= "110000101100";
          WHEN  37 => goldSin <= "000110001001";
                      goldCos <= "110001001110";
          WHEN  38 => goldSin <= "000111100011";
                      goldCos <= "110001111001";
          WHEN  39 => goldSin <= "001000111010";
                      goldCos <= "110010101101";
          WHEN  40 => goldSin <= "001010001010";
                      goldCos <= "110011101001";
          WHEN  41 => goldSin <= "001011010101";
                      goldCos <= "110100101100";
          WHEN  42 => goldSin <= "001100011000";
                      goldCos <= "110101110111";
          WHEN  43 => goldSin <= "001101010100";
                      goldCos <= "110111001000";
          WHEN  44 => goldSin <= "001110000111";
                      goldCos <= "111000011110";
          WHEN  45 => goldSin <= "001110110010";
                      goldCos <= "111001111001";
          WHEN  46 => goldSin <= "001111010100";
                      goldCos <= "111011011000";
          WHEN  47 => goldSin <= "001111101100";
                      goldCos <= "111100111001";
          WHEN  48 => goldSin <= "001111111011";
                      goldCos <= "111110011100";
          WHEN  49 => goldSin <= "010000000000";
                      goldCos <= "000000000001";
          WHEN  50 => goldSin <= "001111111011";
                      goldCos <= "000001100101";
          WHEN  51 => goldSin <= "001111101100";
                      goldCos <= "000011001001";
          WHEN  52 => goldSin <= "001111010100";
                      goldCos <= "000100101010";
          WHEN  53 => goldSin <= "001110110010";
                      goldCos <= "000110001001";
          WHEN  54 => goldSin <= "001110000111";
                      goldCos <= "000111100011";
          WHEN  55 => goldSin <= "001101010011";
                      goldCos <= "001000111010";
          WHEN  56 => goldSin <= "001100010111";
                      goldCos <= "001010001010";
          WHEN  57 => goldSin <= "001011010100";
                      goldCos <= "001011010101";
          WHEN  58 => goldSin <= "001010001001";
                      goldCos <= "001100011000";
          WHEN  59 => goldSin <= "001000111000";
                      goldCos <= "001101010100";
          WHEN  60 => goldSin <= "000111100010";
                      goldCos <= "001110000111";
          WHEN  61 => goldSin <= "000110000111";
                      goldCos <= "001110110010";
          WHEN  62 => goldSin <= "000100101000";
                      goldCos <= "001111010100";
          WHEN  63 => goldSin <= "000011000111";
                      goldCos <= "001111101100";
          WHEN  64 => goldSin <= "000001100100";
                      goldCos <= "001111111011";
          WHEN  65 => goldSin <= "111111101100";
                      goldCos <= "010000000000";
          WHEN  66 => goldSin <= "111101110101";
                      goldCos <= "001111110111";
          WHEN  67 => goldSin <= "111100000000";
                      goldCos <= "001111100000";
          WHEN  68 => goldSin <= "111010001111";
                      goldCos <= "001110111011";
          WHEN  69 => goldSin <= "111000100010";
                      goldCos <= "001110001010";
          WHEN  70 => goldSin <= "110110111100";
                      goldCos <= "001101001100";
          WHEN  71 => goldSin <= "110101011110";
                      goldCos <= "001100000011";
          WHEN  72 => goldSin <= "110100001001";
                      goldCos <= "001010101111";
          WHEN  73 => goldSin <= "110010111110";
                      goldCos <= "001001010010";
          WHEN  74 => goldSin <= "110001111111";
                      goldCos <= "000111101101";
          WHEN  75 => goldSin <= "110001001011";
                      goldCos <= "000110000001";
          WHEN  76 => goldSin <= "110000100101";
                      goldCos <= "000100010000";
          WHEN  77 => goldSin <= "110000001100";
                      goldCos <= "000010011100";
          WHEN  78 => goldSin <= "110000000001";
                      goldCos <= "000000100101";
          WHEN  79 => goldSin <= "110000000011";
                      goldCos <= "111110101110";
          WHEN  80 => goldSin <= "110000010100";
                      goldCos <= "111100110111";
          WHEN  81 => goldSin <= "110000110010";
                      goldCos <= "111011000100";
          WHEN  82 => goldSin <= "110001011101";
                      goldCos <= "111001010101";
          WHEN  83 => goldSin <= "110010010101";
                      goldCos <= "110111101100";
          WHEN  84 => goldSin <= "110011011001";
                      goldCos <= "110110001001";
          WHEN  85 => goldSin <= "110100101000";
                      goldCos <= "110100110000";
          WHEN  86 => goldSin <= "110110000001";
                      goldCos <= "110011100000";
          WHEN  87 => goldSin <= "110111100010";
                      goldCos <= "110010011011";
          WHEN  88 => goldSin <= "111001001011";
                      goldCos <= "110001100010";
          WHEN  89 => goldSin <= "111010111010";
                      goldCos <= "110000110101";
          WHEN  90 => goldSin <= "111100101101";
                      goldCos <= "110000010110";
          WHEN  91 => goldSin <= "111110100011";
                      goldCos <= "110000000100";
          WHEN  92 => goldSin <= "000000011010";
                      goldCos <= "110000000000";
          WHEN  93 => goldSin <= "000010010001";
                      goldCos <= "110000001010";
          WHEN  94 => goldSin <= "000100000110";
                      goldCos <= "110000100010";
          WHEN  95 => goldSin <= "000101110111";
                      goldCos <= "110001000111";
          WHEN  96 => goldSin <= "000111100011";
                      goldCos <= "110001111001";
          WHEN  97 => goldSin <= "001001001001";
                      goldCos <= "110010111000";
          WHEN  98 => goldSin <= "001010100111";
                      goldCos <= "110100000001";
          WHEN  99 => goldSin <= "001011111011";
                      goldCos <= "110101010110";
          WHEN 100 => goldSin <= "001101000110";
                      goldCos <= "110110110011";
          WHEN 101 => goldSin <= "001110000100";
                      goldCos <= "111000011000";
          WHEN 102 => goldSin <= "001110110111";
                      goldCos <= "111010000101";
          WHEN 103 => goldSin <= "001111011101";
                      goldCos <= "111011110110";
          WHEN 104 => goldSin <= "001111110101";
                      goldCos <= "111101101011";
          WHEN 105 => goldSin <= "010000000000";
                      goldCos <= "111111100001";
          WHEN 106 => goldSin <= "001111111100";
                      goldCos <= "000001011001";
          WHEN 107 => goldSin <= "001111101011";
                      goldCos <= "000011001111";
          WHEN 108 => goldSin <= "001111001100";
                      goldCos <= "000101000010";
          WHEN 109 => goldSin <= "001110100000";
                      goldCos <= "000110110001";
          WHEN 110 => goldSin <= "001101100111";
                      goldCos <= "001000011010";
          WHEN 111 => goldSin <= "001100100011";
                      goldCos <= "001001111100";
          WHEN 112 => goldSin <= "001011010100";
                      goldCos <= "001011010101";
          WHEN 113 => goldSin <= "001001111010";
                      goldCos <= "001100100100";
          WHEN 114 => goldSin <= "001000011001";
                      goldCos <= "001101101000";
          WHEN 115 => goldSin <= "000110101111";
                      goldCos <= "001110100001";
          WHEN 116 => goldSin <= "000101000000";
                      goldCos <= "001111001101";
          WHEN 117 => goldSin <= "000011001101";
                      goldCos <= "001111101011";
          WHEN 118 => goldSin <= "000001010111";
                      goldCos <= "001111111100";
          WHEN 119 => goldSin <= "111111100000";
                      goldCos <= "001111111111";
          WHEN 120 => goldSin <= "111101010110";
                      goldCos <= "001111110010";
          WHEN 121 => goldSin <= "111011010000";
                      goldCos <= "001111010010";
          WHEN 122 => goldSin <= "111001001111";
                      goldCos <= "001110100000";
          WHEN 123 => goldSin <= "110111010110";
                      goldCos <= "001101011101";
          WHEN 124 => goldSin <= "110101100111";
                      goldCos <= "001100001011";
          WHEN 125 => goldSin <= "110100000101";
                      goldCos <= "001010101010";
          WHEN 126 => goldSin <= "110010110000";
                      goldCos <= "001000111101";
          WHEN 127 => goldSin <= "110001101010";
                      goldCos <= "000111000110";
          WHEN 128 => goldSin <= "110000110101";
                      goldCos <= "000101000110";
          WHEN 129 => goldSin <= "110000010010";
                      goldCos <= "000011000001";
          WHEN 130 => goldSin <= "110000000010";
                      goldCos <= "000000111000";
          WHEN 131 => goldSin <= "110000000011";
                      goldCos <= "111110101110";
          WHEN 132 => goldSin <= "110000011000";
                      goldCos <= "111100100101";
          WHEN 133 => goldSin <= "110000111110";
                      goldCos <= "111010100000";
          WHEN 134 => goldSin <= "110001110110";
                      goldCos <= "111000100010";
          WHEN 135 => goldSin <= "110010111111";
                      goldCos <= "110110101101";
          WHEN 136 => goldSin <= "110100010111";
                      goldCos <= "110101000010";
          WHEN 137 => goldSin <= "110101111100";
                      goldCos <= "110011100100";
          WHEN 138 => goldSin <= "110111101101";
                      goldCos <= "110010010101";
          WHEN 139 => goldSin <= "111001101000";
                      goldCos <= "110001010101";
          WHEN 140 => goldSin <= "111011101010";
                      goldCos <= "110000100111";
          WHEN 141 => goldSin <= "111101110001";
                      goldCos <= "110000001010";
          WHEN 142 => goldSin <= "111111111011";
                      goldCos <= "110000000000";
          WHEN 143 => goldSin <= "000010000100";
                      goldCos <= "110000001001";
          WHEN 144 => goldSin <= "000100001100";
                      goldCos <= "110000100100";
          WHEN 145 => goldSin <= "000110001110";
                      goldCos <= "110001010001";
          WHEN 146 => goldSin <= "001000001010";
                      goldCos <= "110010001111";
          WHEN 147 => goldSin <= "001001111100";
                      goldCos <= "110011011101";
          WHEN 148 => goldSin <= "001011100010";
                      goldCos <= "110100111010";
          WHEN 149 => goldSin <= "001100111011";
                      goldCos <= "110110100100";
          WHEN 150 => goldSin <= "001110000100";
                      goldCos <= "111000011000";
          WHEN 151 => goldSin <= "001110111110";
                      goldCos <= "111010010110";
          WHEN 152 => goldSin <= "001111100110";
                      goldCos <= "111100011010";
          WHEN 153 => goldSin <= "001111111100";
                      goldCos <= "111110100011";
          WHEN 154 => goldSin <= "001111111111";
                      goldCos <= "000000101101";
          WHEN 155 => goldSin <= "001111110000";
                      goldCos <= "000010110110";
          WHEN 156 => goldSin <= "001111001110";
                      goldCos <= "000100111100";
          WHEN 157 => goldSin <= "001110011011";
                      goldCos <= "000110111100";
          WHEN 158 => goldSin <= "001101010110";
                      goldCos <= "001000110100";
          WHEN 159 => goldSin <= "001100000011";
                      goldCos <= "001010100010";
          WHEN 160 => goldSin <= "001010100001";
                      goldCos <= "001100000100";
          WHEN 161 => goldSin <= "001000110011";
                      goldCos <= "001101010111";
          WHEN 162 => goldSin <= "000110111011";
                      goldCos <= "001110011011";
          WHEN 163 => goldSin <= "000100111010";
                      goldCos <= "001111001111";
          WHEN 164 => goldSin <= "000010110100";
                      goldCos <= "001111110000";
          WHEN 165 => goldSin <= "000000101011";
                      goldCos <= "001111111111";
          WHEN 166 => goldSin <= "111110100001";
                      goldCos <= "001111111100";
          WHEN 167 => goldSin <= "111100011001";
                      goldCos <= "001111100110";
          WHEN 168 => goldSin <= "111010000011";
                      goldCos <= "001110110110";
          WHEN 169 => goldSin <= "110111110110";
                      goldCos <= "001101110001";
          WHEN 170 => goldSin <= "110101110110";
                      goldCos <= "001100010111";
          WHEN 171 => goldSin <= "110100000101";
                      goldCos <= "001010101010";
          WHEN 172 => goldSin <= "110010100101";
                      goldCos <= "001000101110";
          WHEN 173 => goldSin <= "110001011010";
                      goldCos <= "000110100100";
          WHEN 174 => goldSin <= "110000100101";
                      goldCos <= "000100010000";
          WHEN 175 => goldSin <= "110000000111";
                      goldCos <= "000001110110";
          WHEN 176 => goldSin <= "110000000001";
                      goldCos <= "111111011010";
          WHEN 177 => goldSin <= "110000010011";
                      goldCos <= "111100111110";
          WHEN 178 => goldSin <= "110000111100";
                      goldCos <= "111010100110";
          WHEN 179 => goldSin <= "110001111100";
                      goldCos <= "111000010111";
          WHEN 180 => goldSin <= "110011010010";
                      goldCos <= "110110010011";
          WHEN 181 => goldSin <= "110100111010";
                      goldCos <= "110100011110";
          WHEN 182 => goldSin <= "110110110011";
                      goldCos <= "110010111010";
          WHEN 183 => goldSin <= "111000111010";
                      goldCos <= "110001101010";
          WHEN 184 => goldSin <= "111011001011";
                      goldCos <= "110000110000";
          WHEN 185 => goldSin <= "111101100100";
                      goldCos <= "110000001100";
          WHEN 186 => goldSin <= "000000000001";
                      goldCos <= "110000000000";
          WHEN 187 => goldSin <= "000010011101";
                      goldCos <= "110000001100";
          WHEN 188 => goldSin <= "000100110110";
                      goldCos <= "110000110000";
          WHEN 189 => goldSin <= "000111000111";
                      goldCos <= "110001101011";
          WHEN 190 => goldSin <= "001001001110";
                      goldCos <= "110010111011";
          WHEN 191 => goldSin <= "001011000111";
                      goldCos <= "110100011111";
          WHEN 192 => goldSin <= "001100101111";
                      goldCos <= "110110010101";
          WHEN 193 => goldSin <= "001110000100";
                      goldCos <= "111000011000";
          WHEN 194 => goldSin <= "001111000100";
                      goldCos <= "111010101000";
          WHEN 195 => goldSin <= "001111101110";
                      goldCos <= "111100111111";
          WHEN 196 => goldSin <= "001111111111";
                      goldCos <= "111111011011";
          WHEN 197 => goldSin <= "001111111001";
                      goldCos <= "000001111000";
          WHEN 198 => goldSin <= "001111011011";
                      goldCos <= "000100010010";
          WHEN 199 => goldSin <= "001110100101";
                      goldCos <= "000110100101";
          WHEN 200 => goldSin <= "001101011010";
                      goldCos <= "001000101111";
          WHEN 201 => goldSin <= "001011111010";
                      goldCos <= "001010101100";
          WHEN 202 => goldSin <= "001010001001";
                      goldCos <= "001100011000";
          WHEN 203 => goldSin <= "001000001000";
                      goldCos <= "001101110010";
          WHEN 204 => goldSin <= "000101111011";
                      goldCos <= "001110110111";
          WHEN 205 => goldSin <= "000011100110";
                      goldCos <= "001111100110";
          WHEN 206 => goldSin <= "000001001011";
                      goldCos <= "001111111101";
          WHEN 207 => goldSin <= "111110101110";
                      goldCos <= "001111111101";
          WHEN 208 => goldSin <= "111100010011";
                      goldCos <= "001111100100";
          WHEN 209 => goldSin <= "111001111101";
                      goldCos <= "001110110100";
          WHEN 210 => goldSin <= "110111100001";
                      goldCos <= "001101100100";
          WHEN 211 => goldSin <= "110101010100";
                      goldCos <= "001011111010";
          WHEN 212 => goldSin <= "110011011100";
                      goldCos <= "001001111010";
          WHEN 213 => goldSin <= "110001111100";
                      goldCos <= "000111101000";
          WHEN 214 => goldSin <= "110000110101";
                      goldCos <= "000101000110";
          WHEN 215 => goldSin <= "110000001100";
                      goldCos <= "000010011100";
          WHEN 216 => goldSin <= "110000000000";
                      goldCos <= "111111101100";
          WHEN 217 => goldSin <= "110000010011";
                      goldCos <= "111100111110";
          WHEN 218 => goldSin <= "110001000011";
                      goldCos <= "111010010101";
          WHEN 219 => goldSin <= "110010001111";
                      goldCos <= "110111110110";
          WHEN 220 => goldSin <= "110011110101";
                      goldCos <= "110101100111";
          WHEN 221 => goldSin <= "110101110010";
                      goldCos <= "110011101100";
          WHEN 222 => goldSin <= "111000000010";
                      goldCos <= "110010001000";
          WHEN 223 => goldSin <= "111010100010";
                      goldCos <= "110000111110";
          WHEN 224 => goldSin <= "111101001100";
                      goldCos <= "110000010000";
          WHEN 225 => goldSin <= "111111111011";
                      goldCos <= "110000000000";
          WHEN 226 => goldSin <= "000010101010";
                      goldCos <= "110000001110";
          WHEN 227 => goldSin <= "000101010100";
                      goldCos <= "110000111010";
          WHEN 228 => goldSin <= "000111110100";
                      goldCos <= "110010000010";
          WHEN 229 => goldSin <= "001010000101";
                      goldCos <= "110011100101";
          WHEN 230 => goldSin <= "001100000100";
                      goldCos <= "110101011111";
          WHEN 231 => goldSin <= "001101101011";
                      goldCos <= "110111101101";
          WHEN 232 => goldSin <= "001110111001";
                      goldCos <= "111010001010";
          WHEN 233 => goldSin <= "001111101011";
                      goldCos <= "111100110011";
          WHEN 234 => goldSin <= "010000000000";
                      goldCos <= "111111100001";
          WHEN 235 => goldSin <= "001111110110";
                      goldCos <= "000010010001";
          WHEN 236 => goldSin <= "001111001110";
                      goldCos <= "000100111100";
          WHEN 237 => goldSin <= "001110001010";
                      goldCos <= "000111011110";
          WHEN 238 => goldSin <= "001100101011";
                      goldCos <= "001001110010";
          WHEN 239 => goldSin <= "001010110100";
                      goldCos <= "001011110011";
          WHEN 240 => goldSin <= "001000101000";
                      goldCos <= "001101011110";
          WHEN 241 => goldSin <= "000110001101";
                      goldCos <= "001110110000";
          WHEN 242 => goldSin <= "000011100110";
                      goldCos <= "001111100110";
          WHEN 243 => goldSin <= "000000111000";
                      goldCos <= "001111111110";
          WHEN 244 => goldSin <= "111110001000";
                      goldCos <= "001111111001";
          WHEN 245 => goldSin <= "111011011100";
                      goldCos <= "001111010101";
          WHEN 246 => goldSin <= "111000111001";
                      goldCos <= "001110010101";
          WHEN 247 => goldSin <= "110110100010";
                      goldCos <= "001100111010";
          WHEN 248 => goldSin <= "110100010001";
                      goldCos <= "001010111000";
          WHEN 249 => goldSin <= "110010011011";
                      goldCos <= "001000011110";
          WHEN 250 => goldSin <= "110001000100";
                      goldCos <= "000101110000";
          WHEN 251 => goldSin <= "110000010000";
                      goldCos <= "000010110100";
          WHEN 252 => goldSin <= "110000000000";
                      goldCos <= "111111110011";
          WHEN 253 => goldSin <= "110000010101";
                      goldCos <= "111100110001";
          WHEN 254 => goldSin <= "110001001110";
                      goldCos <= "111001110111";
          WHEN 255 => goldSin <= "110010101010";
                      goldCos <= "110111001100";
          WHEN 256 => goldSin <= "110100100100";
                      goldCos <= "110100110100";
          WHEN 257 => goldSin <= "110110111000";
                      goldCos <= "110010110111";
          WHEN 258 => goldSin <= "111001100010";
                      goldCos <= "110001011000";
          WHEN 259 => goldSin <= "111100011010";
                      goldCos <= "110000011010";
          WHEN 260 => goldSin <= "111111011011";
                      goldCos <= "110000000001";
          WHEN 261 => goldSin <= "000010011101";
                      goldCos <= "110000001100";
          WHEN 262 => goldSin <= "000101011010";
                      goldCos <= "110000111100";
          WHEN 263 => goldSin <= "001000001010";
                      goldCos <= "110010001111";
          WHEN 264 => goldSin <= "001010100111";
                      goldCos <= "110100000001";
          WHEN 265 => goldSin <= "001100101100";
                      goldCos <= "110110010000";
          WHEN 266 => goldSin <= "001110010011";
                      goldCos <= "111000110100";
          WHEN 267 => goldSin <= "001111011001";
                      goldCos <= "111011101010";
          WHEN 268 => goldSin <= "001111111100";
                      goldCos <= "111110101001";
          WHEN 269 => goldSin <= "001111111010";
                      goldCos <= "000001101011";
          WHEN 270 => goldSin <= "001111010100";
                      goldCos <= "000100101010";
          WHEN 271 => goldSin <= "001110001010";
                      goldCos <= "000111011110";
          WHEN 272 => goldSin <= "001100011111";
                      goldCos <= "001010000000";
          WHEN 273 => goldSin <= "001010010111";
                      goldCos <= "001100001100";
          WHEN 274 => goldSin <= "000111111000";
                      goldCos <= "001101111011";
          WHEN 275 => goldSin <= "000101000110";
                      goldCos <= "001111001011";
          WHEN 276 => goldSin <= "000010001001";
                      goldCos <= "001111110111";
          WHEN 277 => goldSin <= "111111000111";
                      goldCos <= "001111111110";
          WHEN 278 => goldSin <= "111100000110";
                      goldCos <= "001111100001";
          WHEN 279 => goldSin <= "111001001111";
                      goldCos <= "001110100000";
          WHEN 280 => goldSin <= "110110101000";
                      goldCos <= "001100111101";
          WHEN 281 => goldSin <= "110100010110";
                      goldCos <= "001010111101";
          WHEN 282 => goldSin <= "110010011110";
                      goldCos <= "001000100011";
          WHEN 283 => goldSin <= "110001000000";
                      goldCos <= "000101100100";
          WHEN 284 => goldSin <= "110000001011";
                      goldCos <= "000010010101";
          WHEN 285 => goldSin <= "110000000010";
                      goldCos <= "111111000000";
          WHEN 286 => goldSin <= "110000100101";
                      goldCos <= "111011101110";
          WHEN 287 => goldSin <= "110001110011";
                      goldCos <= "111000101000";
          WHEN 288 => goldSin <= "110011101001";
                      goldCos <= "110101110110";
          WHEN 289 => goldSin <= "110110000001";
                      goldCos <= "110011100000";
          WHEN 290 => goldSin <= "111000110100";
                      goldCos <= "110001101101";
          WHEN 291 => goldSin <= "111011111100";
                      goldCos <= "110000100010";
          WHEN 292 => goldSin <= "111111001111";
                      goldCos <= "110000000001";
          WHEN 293 => goldSin <= "000010100011";
                      goldCos <= "110000001101";
          WHEN 294 => goldSin <= "000101110001";
                      goldCos <= "110001000101";
          WHEN 295 => goldSin <= "001000101111";
                      goldCos <= "110010100110";
          WHEN 296 => goldSin <= "001011010101";
                      goldCos <= "110100101100";
          WHEN 297 => goldSin <= "001101011011";
                      goldCos <= "110111010010";
          WHEN 298 => goldSin <= "001110111100";
                      goldCos <= "111010010000";
          WHEN 299 => goldSin <= "001111110011";
                      goldCos <= "111101011110";
          WHEN 300 => goldSin <= "001111111111";
                      goldCos <= "000000110011";
          WHEN 301 => goldSin <= "001111011110";
                      goldCos <= "000100000110";
          WHEN 302 => goldSin <= "001110010010";
                      goldCos <= "000111001101";
          WHEN 303 => goldSin <= "001100011111";
                      goldCos <= "001010000000";
          WHEN 304 => goldSin <= "001010001001";
                      goldCos <= "001100011000";
          WHEN 305 => goldSin <= "000111010111";
                      goldCos <= "001110001101";
          WHEN 306 => goldSin <= "000100010000";
                      goldCos <= "001111011011";
          WHEN 307 => goldSin <= "000000111110";
                      goldCos <= "001111111110";
          WHEN 308 => goldSin <= "111101101001";
                      goldCos <= "001111110101";
          WHEN 309 => goldSin <= "111010011010";
                      goldCos <= "001111000000";
          WHEN 310 => goldSin <= "110111011011";
                      goldCos <= "001101100001";
          WHEN 311 => goldSin <= "110100110100";
                      goldCos <= "001011011100";
          WHEN 312 => goldSin <= "110010101100";
                      goldCos <= "001000111000";
          WHEN 313 => goldSin <= "110001001001";
                      goldCos <= "000101111011";
          WHEN 314 => goldSin <= "110000001111";
                      goldCos <= "000010101110";
          WHEN 315 => goldSin <= "110000000001";
                      goldCos <= "111111011010";
          WHEN 316 => goldSin <= "110000011111";
                      goldCos <= "111100000110";
          WHEN 317 => goldSin <= "110001101000";
                      goldCos <= "111000111110";
          WHEN 318 => goldSin <= "110011011001";
                      goldCos <= "110110001001";
          WHEN 319 => goldSin <= "110101101101";
                      goldCos <= "110011110000";
          WHEN 320 => goldSin <= "111000011110";
                      goldCos <= "110001111001";
          WHEN 321 => goldSin <= "111011100100";
                      goldCos <= "110000101000";
          WHEN 322 => goldSin <= "111110110101";
                      goldCos <= "110000000011";
          WHEN 323 => goldSin <= "000010001011";
                      goldCos <= "110000001001";
          WHEN 324 => goldSin <= "000101011010";
                      goldCos <= "110000111100";
          WHEN 325 => goldSin <= "001000011010";
                      goldCos <= "110010011001";
          WHEN 326 => goldSin <= "001011000011";
                      goldCos <= "110100011011";
          WHEN 327 => goldSin <= "001101001101";
                      goldCos <= "110110111101";
          WHEN 328 => goldSin <= "001110110010";
                      goldCos <= "111001111001";
          WHEN 329 => goldSin <= "001111101111";
                      goldCos <= "111101000101";
          WHEN 330 => goldSin <= "010000000000";
                      goldCos <= "000000011010";
          WHEN 331 => goldSin <= "001111100100";
                      goldCos <= "000011101101";
          WHEN 332 => goldSin <= "001110011101";
                      goldCos <= "000110110111";
          WHEN 333 => goldSin <= "001100101110";
                      goldCos <= "001001101101";
          WHEN 334 => goldSin <= "001010011100";
                      goldCos <= "001100001000";
          WHEN 335 => goldSin <= "000111101101";
                      goldCos <= "001110000001";
          WHEN 336 => goldSin <= "000100101000";
                      goldCos <= "001111010100";
          WHEN 337 => goldSin <= "000001010111";
                      goldCos <= "001111111100";
          WHEN 338 => goldSin <= "111110000010";
                      goldCos <= "001111111000";
          WHEN 339 => goldSin <= "111010110010";
                      goldCos <= "001111001000";
          WHEN 340 => goldSin <= "110111110001";
                      goldCos <= "001101101110";
          WHEN 341 => goldSin <= "110101000110";
                      goldCos <= "001011101110";
          WHEN 342 => goldSin <= "110010111010";
                      goldCos <= "001001001101";
          WHEN 343 => goldSin <= "110001010011";
                      goldCos <= "000110010011";
          WHEN 344 => goldSin <= "110000010100";
                      goldCos <= "000011000111";
          WHEN 345 => goldSin <= "110000000000";
                      goldCos <= "111111110011";
          WHEN 346 => goldSin <= "110000011001";
                      goldCos <= "111100011111";
          WHEN 347 => goldSin <= "110001011101";
                      goldCos <= "111001010101";
          WHEN 348 => goldSin <= "110011001010";
                      goldCos <= "110110011101";
          WHEN 349 => goldSin <= "110101011010";
                      goldCos <= "110100000000";
          WHEN 350 => goldSin <= "111000001000";
                      goldCos <= "110010000101";
          WHEN 351 => goldSin <= "111011001011";
                      goldCos <= "110000110000";
          WHEN 352 => goldSin <= "111110011100";
                      goldCos <= "110000000101";
          WHEN 353 => goldSin <= "000001110010";
                      goldCos <= "110000000110";
          WHEN 354 => goldSin <= "000101000010";
                      goldCos <= "110000110100";
          WHEN 355 => goldSin <= "001000000100";
                      goldCos <= "110010001100";
          WHEN 356 => goldSin <= "001010110000";
                      goldCos <= "110100001010";
          WHEN 357 => goldSin <= "001100111110";
                      goldCos <= "110110101001";
          WHEN 358 => goldSin <= "001110101000";
                      goldCos <= "111001100010";
          WHEN 359 => goldSin <= "001111101010";
                      goldCos <= "111100101101";
          WHEN 360 => goldSin <= "010000000000";
                      goldCos <= "000000000001";
          WHEN 361 => goldSin <= "001111101010";
                      goldCos <= "000011010101";
          WHEN 362 => goldSin <= "001110101000";
                      goldCos <= "000110100000";
          WHEN 363 => goldSin <= "001100111101";
                      goldCos <= "001001011000";
          WHEN 364 => goldSin <= "001010101111";
                      goldCos <= "001011110111";
          WHEN 365 => goldSin <= "001000000011";
                      goldCos <= "001101110101";
          WHEN 366 => goldSin <= "000101000000";
                      goldCos <= "001111001101";
          WHEN 367 => goldSin <= "000001110000";
                      goldCos <= "001111111010";
          WHEN 368 => goldSin <= "111110011011";
                      goldCos <= "001111111011";
          WHEN 369 => goldSin <= "111011001010";
                      goldCos <= "001111010000";
          WHEN 370 => goldSin <= "111000000111";
                      goldCos <= "001101111011";
          WHEN 371 => goldSin <= "110101011001";
                      goldCos <= "001011111111";
          WHEN 372 => goldSin <= "110011001001";
                      goldCos <= "001001100001";
          WHEN 373 => goldSin <= "110001011101";
                      goldCos <= "000110101010";
          WHEN 374 => goldSin <= "110000011001";
                      goldCos <= "000011100000";
          WHEN 375 => goldSin <= "110000000000";
                      goldCos <= "000000001100";
          WHEN 376 => goldSin <= "110000010100";
                      goldCos <= "111100110111";
          WHEN 377 => goldSin <= "110001010011";
                      goldCos <= "111001101100";
          WHEN 378 => goldSin <= "110010111011";
                      goldCos <= "110110110010";
          WHEN 379 => goldSin <= "110101001000";
                      goldCos <= "110100010001";
          WHEN 380 => goldSin <= "110111110010";
                      goldCos <= "110010010001";
          WHEN 381 => goldSin <= "111010110100";
                      goldCos <= "110000110111";
          WHEN 382 => goldSin <= "111110000011";
                      goldCos <= "110000001000";
          WHEN 383 => goldSin <= "000001011001";
                      goldCos <= "110000000100";
          WHEN 384 => goldSin <= "000100101010";
                      goldCos <= "110000101100";
          WHEN 385 => goldSin <= "000111101110";
                      goldCos <= "110001111111";
          WHEN 386 => goldSin <= "001010011101";
                      goldCos <= "110011111001";
          WHEN 387 => goldSin <= "001100101111";
                      goldCos <= "110110010101";
          WHEN 388 => goldSin <= "001110011110";
                      goldCos <= "111001001011";
          WHEN 389 => goldSin <= "001111100100";
                      goldCos <= "111100010100";
          WHEN 390 => goldSin <= "010000000000";
                      goldCos <= "111111101000";
          WHEN 391 => goldSin <= "001111101111";
                      goldCos <= "000010111100";
          WHEN 392 => goldSin <= "001110110010";
                      goldCos <= "000110001001";
          WHEN 393 => goldSin <= "001101001100";
                      goldCos <= "001001000100";
          WHEN 394 => goldSin <= "001011000010";
                      goldCos <= "001011100110";
          WHEN 395 => goldSin <= "001000011001";
                      goldCos <= "001101101000";
          WHEN 396 => goldSin <= "000101011000";
                      goldCos <= "001111000100";
          WHEN 397 => goldSin <= "000010001001";
                      goldCos <= "001111110111";
          WHEN 398 => goldSin <= "111110110100";
                      goldCos <= "001111111101";
          WHEN 399 => goldSin <= "111011100010";
                      goldCos <= "001111010111";
          WHEN 400 => goldSin <= "111000011101";
                      goldCos <= "001110000111";
          WHEN 401 => goldSin <= "110101101100";
                      goldCos <= "001100001111";
          WHEN 402 => goldSin <= "110011011000";
                      goldCos <= "001001110101";
          WHEN 403 => goldSin <= "110001100111";
                      goldCos <= "000111000000";
          WHEN 404 => goldSin <= "110000011110";
                      goldCos <= "000011111000";
          WHEN 405 => goldSin <= "110000000001";
                      goldCos <= "000000100101";
          WHEN 406 => goldSin <= "110000001111";
                      goldCos <= "111101010000";
          WHEN 407 => goldSin <= "110001001010";
                      goldCos <= "111010000011";
          WHEN 408 => goldSin <= "110010101101";
                      goldCos <= "110111000110";
          WHEN 409 => goldSin <= "110100110101";
                      goldCos <= "110100100011";
          WHEN 410 => goldSin <= "110111011101";
                      goldCos <= "110010011110";
          WHEN 411 => goldSin <= "111010011100";
                      goldCos <= "110001000000";
          WHEN 412 => goldSin <= "111101101011";
                      goldCos <= "110000001011";
          WHEN 413 => goldSin <= "000001000000";
                      goldCos <= "110000000010";
          WHEN 414 => goldSin <= "000100010010";
                      goldCos <= "110000100101";
          WHEN 415 => goldSin <= "000111011000";
                      goldCos <= "110001110011";
          WHEN 416 => goldSin <= "001010001010";
                      goldCos <= "110011101001";
          WHEN 417 => goldSin <= "001100100000";
                      goldCos <= "110110000001";
          WHEN 418 => goldSin <= "001110010011";
                      goldCos <= "111000110100";
          WHEN 419 => goldSin <= "001111011110";
                      goldCos <= "111011111100";
          WHEN 420 => goldSin <= "001111111111";
                      goldCos <= "111111001111";
          WHEN 421 => goldSin <= "001111110011";
                      goldCos <= "000010100011";
          WHEN 422 => goldSin <= "001110111011";
                      goldCos <= "000101110001";
          WHEN 423 => goldSin <= "001101011010";
                      goldCos <= "001000101111";
          WHEN 424 => goldSin <= "001011010100";
                      goldCos <= "001011010101";
          WHEN 425 => goldSin <= "001000101110";
                      goldCos <= "001101011011";
          WHEN 426 => goldSin <= "000101110000";
                      goldCos <= "001110111100";
          WHEN 427 => goldSin <= "000010100010";
                      goldCos <= "001111110011";
          WHEN 428 => goldSin <= "111111001101";
                      goldCos <= "001111111111";
          WHEN 429 => goldSin <= "111011111010";
                      goldCos <= "001111011110";
          WHEN 430 => goldSin <= "111000110011";
                      goldCos <= "001110010010";
          WHEN 431 => goldSin <= "110110000000";
                      goldCos <= "001100011111";
          WHEN 432 => goldSin <= "110011101000";
                      goldCos <= "001010001001";
          WHEN 433 => goldSin <= "110001110011";
                      goldCos <= "000111010111";
          WHEN 434 => goldSin <= "110000100101";
                      goldCos <= "000100010000";
          WHEN 435 => goldSin <= "110000000010";
                      goldCos <= "000000111110";
          WHEN 436 => goldSin <= "110000001011";
                      goldCos <= "111101101001";
          WHEN 437 => goldSin <= "110001000000";
                      goldCos <= "111010011010";
          WHEN 438 => goldSin <= "110010011111";
                      goldCos <= "110111011011";
          WHEN 439 => goldSin <= "110100100100";
                      goldCos <= "110100110100";
          WHEN 440 => goldSin <= "110111001000";
                      goldCos <= "110010101100";
          WHEN 441 => goldSin <= "111010000101";
                      goldCos <= "110001001001";
          WHEN 442 => goldSin <= "111101010010";
                      goldCos <= "110000001111";
          WHEN 443 => goldSin <= "000000100110";
                      goldCos <= "110000000001";
          WHEN 444 => goldSin <= "000011111010";
                      goldCos <= "110000011111";
          WHEN 445 => goldSin <= "000111000010";
                      goldCos <= "110001101000";
          WHEN 446 => goldSin <= "001001110111";
                      goldCos <= "110011011001";
          WHEN 447 => goldSin <= "001100010000";
                      goldCos <= "110101101101";
          WHEN 448 => goldSin <= "001110000111";
                      goldCos <= "111000011110";
          WHEN 449 => goldSin <= "001111011000";
                      goldCos <= "111011100100";
          WHEN 450 => goldSin <= "001111111101";
                      goldCos <= "111110110101";
          WHEN 451 => goldSin <= "001111110111";
                      goldCos <= "000010001011";
          WHEN 452 => goldSin <= "001111000100";
                      goldCos <= "000101011010";
          WHEN 453 => goldSin <= "001101100111";
                      goldCos <= "001000011010";
          WHEN 454 => goldSin <= "001011100101";
                      goldCos <= "001011000011";
          WHEN 455 => goldSin <= "001001000011";
                      goldCos <= "001101001101";
          WHEN 456 => goldSin <= "000110000111";
                      goldCos <= "001110110010";
          WHEN 457 => goldSin <= "000010111011";
                      goldCos <= "001111101111";
          WHEN 458 => goldSin <= "111111100110";
                      goldCos <= "010000000000";
          WHEN 459 => goldSin <= "111100010011";
                      goldCos <= "001111100100";
          WHEN 460 => goldSin <= "111001001001";
                      goldCos <= "001110011101";
          WHEN 461 => goldSin <= "110110010011";
                      goldCos <= "001100101110";
          WHEN 462 => goldSin <= "110011111000";
                      goldCos <= "001010011100";
          WHEN 463 => goldSin <= "110001111111";
                      goldCos <= "000111101101";
          WHEN 464 => goldSin <= "110000101100";
                      goldCos <= "000100101000";
          WHEN 465 => goldSin <= "110000000100";
                      goldCos <= "000001010111";
          WHEN 466 => goldSin <= "110000001000";
                      goldCos <= "111110000010";
          WHEN 467 => goldSin <= "110000111000";
                      goldCos <= "111010110010";
          WHEN 468 => goldSin <= "110010010010";
                      goldCos <= "110111110001";
          WHEN 469 => goldSin <= "110100010010";
                      goldCos <= "110101000110";
          WHEN 470 => goldSin <= "110110110011";
                      goldCos <= "110010111010";
          WHEN 471 => goldSin <= "111001101101";
                      goldCos <= "110001010011";
          WHEN 472 => goldSin <= "111100111001";
                      goldCos <= "110000010100";
          WHEN 473 => goldSin <= "000000001101";
                      goldCos <= "110000000000";
          WHEN 474 => goldSin <= "000011100001";
                      goldCos <= "110000011001";
          WHEN 475 => goldSin <= "000110101011";
                      goldCos <= "110001011101";
          WHEN 476 => goldSin <= "001001100011";
                      goldCos <= "110011001010";
          WHEN 477 => goldSin <= "001100000000";
                      goldCos <= "110101011010";
          WHEN 478 => goldSin <= "001101111011";
                      goldCos <= "111000001000";
          WHEN 479 => goldSin <= "001111010000";
                      goldCos <= "111011001011";
          WHEN 480 => goldSin <= "001111111011";
                      goldCos <= "111110011100";
          WHEN 481 => goldSin <= "001111111010";
                      goldCos <= "000001110010";
          WHEN 482 => goldSin <= "001111001100";
                      goldCos <= "000101000010";
          WHEN 483 => goldSin <= "001101110100";
                      goldCos <= "001000000100";
          WHEN 484 => goldSin <= "001011110110";
                      goldCos <= "001010110000";
          WHEN 485 => goldSin <= "001001010111";
                      goldCos <= "001100111110";
          WHEN 486 => goldSin <= "000110011110";
                      goldCos <= "001110101000";
          WHEN 487 => goldSin <= "000011010011";
                      goldCos <= "001111101010";
          WHEN 488 => goldSin <= "111111111111";
                      goldCos <= "010000000000";
          WHEN 489 => goldSin <= "111100101011";
                      goldCos <= "001111101010";
          WHEN 490 => goldSin <= "111001100000";
                      goldCos <= "001110101000";
          WHEN 491 => goldSin <= "110110101000";
                      goldCos <= "001100111101";
          WHEN 492 => goldSin <= "110100001001";
                      goldCos <= "001010101111";
          WHEN 493 => goldSin <= "110010001011";
                      goldCos <= "001000000011";
          WHEN 494 => goldSin <= "110000110011";
                      goldCos <= "000101000000";
          WHEN 495 => goldSin <= "110000000110";
                      goldCos <= "000001110000";
          WHEN 496 => goldSin <= "110000000101";
                      goldCos <= "111110011011";
          WHEN 497 => goldSin <= "110000110000";
                      goldCos <= "111011001010";
          WHEN 498 => goldSin <= "110010000101";
                      goldCos <= "111000000111";
          WHEN 499 => goldSin <= "110100000001";
                      goldCos <= "110101011001";
          WHEN 500 => goldSin <= "110110011111";
                      goldCos <= "110011001001";
          WHEN 501 => goldSin <= "111001010110";
                      goldCos <= "110001011101";
          WHEN 502 => goldSin <= "111100100000";
                      goldCos <= "110000011001";
          WHEN 503 => goldSin <= "111111110100";
                      goldCos <= "110000000000";
          WHEN 504 => goldSin <= "000011001001";
                      goldCos <= "110000010100";
          WHEN 505 => goldSin <= "000110010100";
                      goldCos <= "110001010011";
          WHEN 506 => goldSin <= "001001001110";
                      goldCos <= "110010111011";
          WHEN 507 => goldSin <= "001011101111";
                      goldCos <= "110101001000";
          WHEN 508 => goldSin <= "001101101111";
                      goldCos <= "110111110010";
          WHEN 509 => goldSin <= "001111001001";
                      goldCos <= "111010110100";
       WHEN OTHERS => goldSin <= (others=>'0');
                      goldCos <= (others=>'0');
        END CASE; 
    END PROCESS; 
END ARCHITECTURE rtl; 



