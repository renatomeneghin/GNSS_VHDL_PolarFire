LIBRARY IEEE; 
  USE IEEE.std_logic_1164.all; 
  USE IEEE.numeric_std.all; 

ENTITY COREDDS_C0_COREDDS_C0_0_dds_qrtr_sin IS 
  PORT ( 
    index : IN std_logic_vector(8 DOWNTO 0); 
    sine : OUT std_logic_vector(11 DOWNTO 0)); 

    attribute syn_noclockbuf: Boolean;                    --03/09/17 
    attribute syn_noclockbuf of index : signal is true;   --03/09/17 
    attribute syn_noclockbuf of sine  : signal is true;   --03/09/17 
END ENTITY COREDDS_C0_COREDDS_C0_0_dds_qrtr_sin; 

ARCHITECTURE rtl OF COREDDS_C0_COREDDS_C0_0_dds_qrtr_sin IS 
  SIGNAL A_int : integer; 
BEGIN 
  A_int <= to_integer(unsigned(index)); 
  PROCESS (A_int) 
    VARIABLE wave : std_logic_vector(11 DOWNTO 0); 
  BEGIN 
    CASE A_int IS      -- synopsys parallel_case     
      WHEN    0 => wave := "000000000001"; --          1 
      WHEN    1 => wave := "000000000010"; --          2 
      WHEN    2 => wave := "000000000100"; --          4 
      WHEN    3 => wave := "000000000101"; --          5 
      WHEN    4 => wave := "000000000111"; --          7 
      WHEN    5 => wave := "000000001001"; --          9 
      WHEN    6 => wave := "000000001010"; --         10 
      WHEN    7 => wave := "000000001100"; --         12 
      WHEN    8 => wave := "000000001101"; --         13 
      WHEN    9 => wave := "000000001111"; --         15 
      WHEN   10 => wave := "000000010000"; --         16 
      WHEN   11 => wave := "000000010010"; --         18 
      WHEN   12 => wave := "000000010100"; --         20 
      WHEN   13 => wave := "000000010101"; --         21 
      WHEN   14 => wave := "000000010111"; --         23 
      WHEN   15 => wave := "000000011000"; --         24 
      WHEN   16 => wave := "000000011010"; --         26 
      WHEN   17 => wave := "000000011011"; --         27 
      WHEN   18 => wave := "000000011101"; --         29 
      WHEN   19 => wave := "000000011111"; --         31 
      WHEN   20 => wave := "000000100000"; --         32 
      WHEN   21 => wave := "000000100010"; --         34 
      WHEN   22 => wave := "000000100011"; --         35 
      WHEN   23 => wave := "000000100101"; --         37 
      WHEN   24 => wave := "000000100110"; --         38 
      WHEN   25 => wave := "000000101000"; --         40 
      WHEN   26 => wave := "000000101010"; --         42 
      WHEN   27 => wave := "000000101011"; --         43 
      WHEN   28 => wave := "000000101101"; --         45 
      WHEN   29 => wave := "000000101110"; --         46 
      WHEN   30 => wave := "000000110000"; --         48 
      WHEN   31 => wave := "000000110001"; --         49 
      WHEN   32 => wave := "000000110011"; --         51 
      WHEN   33 => wave := "000000110101"; --         53 
      WHEN   34 => wave := "000000110110"; --         54 
      WHEN   35 => wave := "000000111000"; --         56 
      WHEN   36 => wave := "000000111001"; --         57 
      WHEN   37 => wave := "000000111011"; --         59 
      WHEN   38 => wave := "000000111100"; --         60 
      WHEN   39 => wave := "000000111110"; --         62 
      WHEN   40 => wave := "000001000000"; --         64 
      WHEN   41 => wave := "000001000001"; --         65 
      WHEN   42 => wave := "000001000011"; --         67 
      WHEN   43 => wave := "000001000100"; --         68 
      WHEN   44 => wave := "000001000110"; --         70 
      WHEN   45 => wave := "000001000111"; --         71 
      WHEN   46 => wave := "000001001001"; --         73 
      WHEN   47 => wave := "000001001011"; --         75 
      WHEN   48 => wave := "000001001100"; --         76 
      WHEN   49 => wave := "000001001110"; --         78 
      WHEN   50 => wave := "000001001111"; --         79 
      WHEN   51 => wave := "000001010001"; --         81 
      WHEN   52 => wave := "000001010010"; --         82 
      WHEN   53 => wave := "000001010100"; --         84 
      WHEN   54 => wave := "000001010110"; --         86 
      WHEN   55 => wave := "000001010111"; --         87 
      WHEN   56 => wave := "000001011001"; --         89 
      WHEN   57 => wave := "000001011010"; --         90 
      WHEN   58 => wave := "000001011100"; --         92 
      WHEN   59 => wave := "000001011101"; --         93 
      WHEN   60 => wave := "000001011111"; --         95 
      WHEN   61 => wave := "000001100000"; --         96 
      WHEN   62 => wave := "000001100010"; --         98 
      WHEN   63 => wave := "000001100100"; --        100 
      WHEN   64 => wave := "000001100101"; --        101 
      WHEN   65 => wave := "000001100111"; --        103 
      WHEN   66 => wave := "000001101000"; --        104 
      WHEN   67 => wave := "000001101010"; --        106 
      WHEN   68 => wave := "000001101011"; --        107 
      WHEN   69 => wave := "000001101101"; --        109 
      WHEN   70 => wave := "000001101111"; --        111 
      WHEN   71 => wave := "000001110000"; --        112 
      WHEN   72 => wave := "000001110010"; --        114 
      WHEN   73 => wave := "000001110011"; --        115 
      WHEN   74 => wave := "000001110101"; --        117 
      WHEN   75 => wave := "000001110110"; --        118 
      WHEN   76 => wave := "000001111000"; --        120 
      WHEN   77 => wave := "000001111001"; --        121 
      WHEN   78 => wave := "000001111011"; --        123 
      WHEN   79 => wave := "000001111101"; --        125 
      WHEN   80 => wave := "000001111110"; --        126 
      WHEN   81 => wave := "000010000000"; --        128 
      WHEN   82 => wave := "000010000001"; --        129 
      WHEN   83 => wave := "000010000011"; --        131 
      WHEN   84 => wave := "000010000100"; --        132 
      WHEN   85 => wave := "000010000110"; --        134 
      WHEN   86 => wave := "000010000111"; --        135 
      WHEN   87 => wave := "000010001001"; --        137 
      WHEN   88 => wave := "000010001011"; --        139 
      WHEN   89 => wave := "000010001100"; --        140 
      WHEN   90 => wave := "000010001110"; --        142 
      WHEN   91 => wave := "000010001111"; --        143 
      WHEN   92 => wave := "000010010001"; --        145 
      WHEN   93 => wave := "000010010010"; --        146 
      WHEN   94 => wave := "000010010100"; --        148 
      WHEN   95 => wave := "000010010101"; --        149 
      WHEN   96 => wave := "000010010111"; --        151 
      WHEN   97 => wave := "000010011001"; --        153 
      WHEN   98 => wave := "000010011010"; --        154 
      WHEN   99 => wave := "000010011100"; --        156 
      WHEN  100 => wave := "000010011101"; --        157 
      WHEN  101 => wave := "000010011111"; --        159 
      WHEN  102 => wave := "000010100000"; --        160 
      WHEN  103 => wave := "000010100010"; --        162 
      WHEN  104 => wave := "000010100011"; --        163 
      WHEN  105 => wave := "000010100101"; --        165 
      WHEN  106 => wave := "000010100111"; --        167 
      WHEN  107 => wave := "000010101000"; --        168 
      WHEN  108 => wave := "000010101010"; --        170 
      WHEN  109 => wave := "000010101011"; --        171 
      WHEN  110 => wave := "000010101101"; --        173 
      WHEN  111 => wave := "000010101110"; --        174 
      WHEN  112 => wave := "000010110000"; --        176 
      WHEN  113 => wave := "000010110001"; --        177 
      WHEN  114 => wave := "000010110011"; --        179 
      WHEN  115 => wave := "000010110100"; --        180 
      WHEN  116 => wave := "000010110110"; --        182 
      WHEN  117 => wave := "000010111000"; --        184 
      WHEN  118 => wave := "000010111001"; --        185 
      WHEN  119 => wave := "000010111011"; --        187 
      WHEN  120 => wave := "000010111100"; --        188 
      WHEN  121 => wave := "000010111110"; --        190 
      WHEN  122 => wave := "000010111111"; --        191 
      WHEN  123 => wave := "000011000001"; --        193 
      WHEN  124 => wave := "000011000010"; --        194 
      WHEN  125 => wave := "000011000100"; --        196 
      WHEN  126 => wave := "000011000101"; --        197 
      WHEN  127 => wave := "000011000111"; --        199 
      WHEN  128 => wave := "000011001001"; --        201 
      WHEN  129 => wave := "000011001010"; --        202 
      WHEN  130 => wave := "000011001100"; --        204 
      WHEN  131 => wave := "000011001101"; --        205 
      WHEN  132 => wave := "000011001111"; --        207 
      WHEN  133 => wave := "000011010000"; --        208 
      WHEN  134 => wave := "000011010010"; --        210 
      WHEN  135 => wave := "000011010011"; --        211 
      WHEN  136 => wave := "000011010101"; --        213 
      WHEN  137 => wave := "000011010110"; --        214 
      WHEN  138 => wave := "000011011000"; --        216 
      WHEN  139 => wave := "000011011001"; --        217 
      WHEN  140 => wave := "000011011011"; --        219 
      WHEN  141 => wave := "000011011101"; --        221 
      WHEN  142 => wave := "000011011110"; --        222 
      WHEN  143 => wave := "000011100000"; --        224 
      WHEN  144 => wave := "000011100001"; --        225 
      WHEN  145 => wave := "000011100011"; --        227 
      WHEN  146 => wave := "000011100100"; --        228 
      WHEN  147 => wave := "000011100110"; --        230 
      WHEN  148 => wave := "000011100111"; --        231 
      WHEN  149 => wave := "000011101001"; --        233 
      WHEN  150 => wave := "000011101010"; --        234 
      WHEN  151 => wave := "000011101100"; --        236 
      WHEN  152 => wave := "000011101101"; --        237 
      WHEN  153 => wave := "000011101111"; --        239 
      WHEN  154 => wave := "000011110000"; --        240 
      WHEN  155 => wave := "000011110010"; --        242 
      WHEN  156 => wave := "000011110011"; --        243 
      WHEN  157 => wave := "000011110101"; --        245 
      WHEN  158 => wave := "000011110111"; --        247 
      WHEN  159 => wave := "000011111000"; --        248 
      WHEN  160 => wave := "000011111010"; --        250 
      WHEN  161 => wave := "000011111011"; --        251 
      WHEN  162 => wave := "000011111101"; --        253 
      WHEN  163 => wave := "000011111110"; --        254 
      WHEN  164 => wave := "000100000000"; --        256 
      WHEN  165 => wave := "000100000001"; --        257 
      WHEN  166 => wave := "000100000011"; --        259 
      WHEN  167 => wave := "000100000100"; --        260 
      WHEN  168 => wave := "000100000110"; --        262 
      WHEN  169 => wave := "000100000111"; --        263 
      WHEN  170 => wave := "000100001001"; --        265 
      WHEN  171 => wave := "000100001010"; --        266 
      WHEN  172 => wave := "000100001100"; --        268 
      WHEN  173 => wave := "000100001101"; --        269 
      WHEN  174 => wave := "000100001111"; --        271 
      WHEN  175 => wave := "000100010000"; --        272 
      WHEN  176 => wave := "000100010010"; --        274 
      WHEN  177 => wave := "000100010011"; --        275 
      WHEN  178 => wave := "000100010101"; --        277 
      WHEN  179 => wave := "000100010110"; --        278 
      WHEN  180 => wave := "000100011000"; --        280 
      WHEN  181 => wave := "000100011001"; --        281 
      WHEN  182 => wave := "000100011011"; --        283 
      WHEN  183 => wave := "000100011100"; --        284 
      WHEN  184 => wave := "000100011110"; --        286 
      WHEN  185 => wave := "000100011111"; --        287 
      WHEN  186 => wave := "000100100001"; --        289 
      WHEN  187 => wave := "000100100010"; --        290 
      WHEN  188 => wave := "000100100100"; --        292 
      WHEN  189 => wave := "000100100101"; --        293 
      WHEN  190 => wave := "000100100111"; --        295 
      WHEN  191 => wave := "000100101000"; --        296 
      WHEN  192 => wave := "000100101010"; --        298 
      WHEN  193 => wave := "000100101100"; --        300 
      WHEN  194 => wave := "000100101101"; --        301 
      WHEN  195 => wave := "000100101111"; --        303 
      WHEN  196 => wave := "000100110000"; --        304 
      WHEN  197 => wave := "000100110010"; --        306 
      WHEN  198 => wave := "000100110011"; --        307 
      WHEN  199 => wave := "000100110101"; --        309 
      WHEN  200 => wave := "000100110110"; --        310 
      WHEN  201 => wave := "000100110111"; --        311 
      WHEN  202 => wave := "000100111001"; --        313 
      WHEN  203 => wave := "000100111010"; --        314 
      WHEN  204 => wave := "000100111100"; --        316 
      WHEN  205 => wave := "000100111101"; --        317 
      WHEN  206 => wave := "000100111111"; --        319 
      WHEN  207 => wave := "000101000000"; --        320 
      WHEN  208 => wave := "000101000010"; --        322 
      WHEN  209 => wave := "000101000011"; --        323 
      WHEN  210 => wave := "000101000101"; --        325 
      WHEN  211 => wave := "000101000110"; --        326 
      WHEN  212 => wave := "000101001000"; --        328 
      WHEN  213 => wave := "000101001001"; --        329 
      WHEN  214 => wave := "000101001011"; --        331 
      WHEN  215 => wave := "000101001100"; --        332 
      WHEN  216 => wave := "000101001110"; --        334 
      WHEN  217 => wave := "000101001111"; --        335 
      WHEN  218 => wave := "000101010001"; --        337 
      WHEN  219 => wave := "000101010010"; --        338 
      WHEN  220 => wave := "000101010100"; --        340 
      WHEN  221 => wave := "000101010101"; --        341 
      WHEN  222 => wave := "000101010111"; --        343 
      WHEN  223 => wave := "000101011000"; --        344 
      WHEN  224 => wave := "000101011010"; --        346 
      WHEN  225 => wave := "000101011011"; --        347 
      WHEN  226 => wave := "000101011101"; --        349 
      WHEN  227 => wave := "000101011110"; --        350 
      WHEN  228 => wave := "000101100000"; --        352 
      WHEN  229 => wave := "000101100001"; --        353 
      WHEN  230 => wave := "000101100011"; --        355 
      WHEN  231 => wave := "000101100100"; --        356 
      WHEN  232 => wave := "000101100110"; --        358 
      WHEN  233 => wave := "000101100111"; --        359 
      WHEN  234 => wave := "000101101000"; --        360 
      WHEN  235 => wave := "000101101010"; --        362 
      WHEN  236 => wave := "000101101011"; --        363 
      WHEN  237 => wave := "000101101101"; --        365 
      WHEN  238 => wave := "000101101110"; --        366 
      WHEN  239 => wave := "000101110000"; --        368 
      WHEN  240 => wave := "000101110001"; --        369 
      WHEN  241 => wave := "000101110011"; --        371 
      WHEN  242 => wave := "000101110100"; --        372 
      WHEN  243 => wave := "000101110110"; --        374 
      WHEN  244 => wave := "000101110111"; --        375 
      WHEN  245 => wave := "000101111001"; --        377 
      WHEN  246 => wave := "000101111010"; --        378 
      WHEN  247 => wave := "000101111011"; --        379 
      WHEN  248 => wave := "000101111101"; --        381 
      WHEN  249 => wave := "000101111110"; --        382 
      WHEN  250 => wave := "000110000000"; --        384 
      WHEN  251 => wave := "000110000001"; --        385 
      WHEN  252 => wave := "000110000011"; --        387 
      WHEN  253 => wave := "000110000100"; --        388 
      WHEN  254 => wave := "000110000110"; --        390 
      WHEN  255 => wave := "000110000111"; --        391 
      WHEN  256 => wave := "000110001001"; --        393 
      WHEN  257 => wave := "000110001010"; --        394 
      WHEN  258 => wave := "000110001011"; --        395 
      WHEN  259 => wave := "000110001101"; --        397 
      WHEN  260 => wave := "000110001110"; --        398 
      WHEN  261 => wave := "000110010000"; --        400 
      WHEN  262 => wave := "000110010001"; --        401 
      WHEN  263 => wave := "000110010011"; --        403 
      WHEN  264 => wave := "000110010100"; --        404 
      WHEN  265 => wave := "000110010110"; --        406 
      WHEN  266 => wave := "000110010111"; --        407 
      WHEN  267 => wave := "000110011000"; --        408 
      WHEN  268 => wave := "000110011010"; --        410 
      WHEN  269 => wave := "000110011011"; --        411 
      WHEN  270 => wave := "000110011101"; --        413 
      WHEN  271 => wave := "000110011110"; --        414 
      WHEN  272 => wave := "000110100000"; --        416 
      WHEN  273 => wave := "000110100001"; --        417 
      WHEN  274 => wave := "000110100011"; --        419 
      WHEN  275 => wave := "000110100100"; --        420 
      WHEN  276 => wave := "000110100101"; --        421 
      WHEN  277 => wave := "000110100111"; --        423 
      WHEN  278 => wave := "000110101000"; --        424 
      WHEN  279 => wave := "000110101010"; --        426 
      WHEN  280 => wave := "000110101011"; --        427 
      WHEN  281 => wave := "000110101101"; --        429 
      WHEN  282 => wave := "000110101110"; --        430 
      WHEN  283 => wave := "000110101111"; --        431 
      WHEN  284 => wave := "000110110001"; --        433 
      WHEN  285 => wave := "000110110010"; --        434 
      WHEN  286 => wave := "000110110100"; --        436 
      WHEN  287 => wave := "000110110101"; --        437 
      WHEN  288 => wave := "000110110111"; --        439 
      WHEN  289 => wave := "000110111000"; --        440 
      WHEN  290 => wave := "000110111001"; --        441 
      WHEN  291 => wave := "000110111011"; --        443 
      WHEN  292 => wave := "000110111100"; --        444 
      WHEN  293 => wave := "000110111110"; --        446 
      WHEN  294 => wave := "000110111111"; --        447 
      WHEN  295 => wave := "000111000000"; --        448 
      WHEN  296 => wave := "000111000010"; --        450 
      WHEN  297 => wave := "000111000011"; --        451 
      WHEN  298 => wave := "000111000101"; --        453 
      WHEN  299 => wave := "000111000110"; --        454 
      WHEN  300 => wave := "000111000111"; --        455 
      WHEN  301 => wave := "000111001001"; --        457 
      WHEN  302 => wave := "000111001010"; --        458 
      WHEN  303 => wave := "000111001100"; --        460 
      WHEN  304 => wave := "000111001101"; --        461 
      WHEN  305 => wave := "000111001111"; --        463 
      WHEN  306 => wave := "000111010000"; --        464 
      WHEN  307 => wave := "000111010001"; --        465 
      WHEN  308 => wave := "000111010011"; --        467 
      WHEN  309 => wave := "000111010100"; --        468 
      WHEN  310 => wave := "000111010101"; --        469 
      WHEN  311 => wave := "000111010111"; --        471 
      WHEN  312 => wave := "000111011000"; --        472 
      WHEN  313 => wave := "000111011010"; --        474 
      WHEN  314 => wave := "000111011011"; --        475 
      WHEN  315 => wave := "000111011100"; --        476 
      WHEN  316 => wave := "000111011110"; --        478 
      WHEN  317 => wave := "000111011111"; --        479 
      WHEN  318 => wave := "000111100001"; --        481 
      WHEN  319 => wave := "000111100010"; --        482 
      WHEN  320 => wave := "000111100011"; --        483 
      WHEN  321 => wave := "000111100101"; --        485 
      WHEN  322 => wave := "000111100110"; --        486 
      WHEN  323 => wave := "000111101000"; --        488 
      WHEN  324 => wave := "000111101001"; --        489 
      WHEN  325 => wave := "000111101010"; --        490 
      WHEN  326 => wave := "000111101100"; --        492 
      WHEN  327 => wave := "000111101101"; --        493 
      WHEN  328 => wave := "000111101110"; --        494 
      WHEN  329 => wave := "000111110000"; --        496 
      WHEN  330 => wave := "000111110001"; --        497 
      WHEN  331 => wave := "000111110011"; --        499 
      WHEN  332 => wave := "000111110100"; --        500 
      WHEN  333 => wave := "000111110101"; --        501 
      WHEN  334 => wave := "000111110111"; --        503 
      WHEN  335 => wave := "000111111000"; --        504 
      WHEN  336 => wave := "000111111001"; --        505 
      WHEN  337 => wave := "000111111011"; --        507 
      WHEN  338 => wave := "000111111100"; --        508 
      WHEN  339 => wave := "000111111110"; --        510 
      WHEN  340 => wave := "000111111111"; --        511 
      WHEN  341 => wave := "001000000000"; --        512 
      WHEN  342 => wave := "001000000010"; --        514 
      WHEN  343 => wave := "001000000011"; --        515 
      WHEN  344 => wave := "001000000100"; --        516 
      WHEN  345 => wave := "001000000110"; --        518 
      WHEN  346 => wave := "001000000111"; --        519 
      WHEN  347 => wave := "001000001000"; --        520 
      WHEN  348 => wave := "001000001010"; --        522 
      WHEN  349 => wave := "001000001011"; --        523 
      WHEN  350 => wave := "001000001100"; --        524 
      WHEN  351 => wave := "001000001110"; --        526 
      WHEN  352 => wave := "001000001111"; --        527 
      WHEN  353 => wave := "001000010000"; --        528 
      WHEN  354 => wave := "001000010010"; --        530 
      WHEN  355 => wave := "001000010011"; --        531 
      WHEN  356 => wave := "001000010100"; --        532 
      WHEN  357 => wave := "001000010110"; --        534 
      WHEN  358 => wave := "001000010111"; --        535 
      WHEN  359 => wave := "001000011001"; --        537 
      WHEN  360 => wave := "001000011010"; --        538 
      WHEN  361 => wave := "001000011011"; --        539 
      WHEN  362 => wave := "001000011101"; --        541 
      WHEN  363 => wave := "001000011110"; --        542 
      WHEN  364 => wave := "001000011111"; --        543 
      WHEN  365 => wave := "001000100001"; --        545 
      WHEN  366 => wave := "001000100010"; --        546 
      WHEN  367 => wave := "001000100011"; --        547 
      WHEN  368 => wave := "001000100101"; --        549 
      WHEN  369 => wave := "001000100110"; --        550 
      WHEN  370 => wave := "001000100111"; --        551 
      WHEN  371 => wave := "001000101000"; --        552 
      WHEN  372 => wave := "001000101010"; --        554 
      WHEN  373 => wave := "001000101011"; --        555 
      WHEN  374 => wave := "001000101100"; --        556 
      WHEN  375 => wave := "001000101110"; --        558 
      WHEN  376 => wave := "001000101111"; --        559 
      WHEN  377 => wave := "001000110000"; --        560 
      WHEN  378 => wave := "001000110010"; --        562 
      WHEN  379 => wave := "001000110011"; --        563 
      WHEN  380 => wave := "001000110100"; --        564 
      WHEN  381 => wave := "001000110110"; --        566 
      WHEN  382 => wave := "001000110111"; --        567 
      WHEN  383 => wave := "001000111000"; --        568 
      WHEN  384 => wave := "001000111010"; --        570 
      WHEN  385 => wave := "001000111011"; --        571 
      WHEN  386 => wave := "001000111100"; --        572 
      WHEN  387 => wave := "001000111101"; --        573 
      WHEN  388 => wave := "001000111111"; --        575 
      WHEN  389 => wave := "001001000000"; --        576 
      WHEN  390 => wave := "001001000001"; --        577 
      WHEN  391 => wave := "001001000011"; --        579 
      WHEN  392 => wave := "001001000100"; --        580 
      WHEN  393 => wave := "001001000101"; --        581 
      WHEN  394 => wave := "001001000111"; --        583 
      WHEN  395 => wave := "001001001000"; --        584 
      WHEN  396 => wave := "001001001001"; --        585 
      WHEN  397 => wave := "001001001010"; --        586 
      WHEN  398 => wave := "001001001100"; --        588 
      WHEN  399 => wave := "001001001101"; --        589 
      WHEN  400 => wave := "001001001110"; --        590 
      WHEN  401 => wave := "001001010000"; --        592 
      WHEN  402 => wave := "001001010001"; --        593 
      WHEN  403 => wave := "001001010010"; --        594 
      WHEN  404 => wave := "001001010011"; --        595 
      WHEN  405 => wave := "001001010101"; --        597 
      WHEN  406 => wave := "001001010110"; --        598 
      WHEN  407 => wave := "001001010111"; --        599 
      WHEN  408 => wave := "001001011000"; --        600 
      WHEN  409 => wave := "001001011010"; --        602 
      WHEN  410 => wave := "001001011011"; --        603 
      WHEN  411 => wave := "001001011100"; --        604 
      WHEN  412 => wave := "001001011110"; --        606 
      WHEN  413 => wave := "001001011111"; --        607 
      WHEN  414 => wave := "001001100000"; --        608 
      WHEN  415 => wave := "001001100001"; --        609 
      WHEN  416 => wave := "001001100011"; --        611 
      WHEN  417 => wave := "001001100100"; --        612 
      WHEN  418 => wave := "001001100101"; --        613 
      WHEN  419 => wave := "001001100110"; --        614 
      WHEN  420 => wave := "001001101000"; --        616 
      WHEN  421 => wave := "001001101001"; --        617 
      WHEN  422 => wave := "001001101010"; --        618 
      WHEN  423 => wave := "001001101011"; --        619 
      WHEN  424 => wave := "001001101101"; --        621 
      WHEN  425 => wave := "001001101110"; --        622 
      WHEN  426 => wave := "001001101111"; --        623 
      WHEN  427 => wave := "001001110000"; --        624 
      WHEN  428 => wave := "001001110010"; --        626 
      WHEN  429 => wave := "001001110011"; --        627 
      WHEN  430 => wave := "001001110100"; --        628 
      WHEN  431 => wave := "001001110101"; --        629 
      WHEN  432 => wave := "001001110111"; --        631 
      WHEN  433 => wave := "001001111000"; --        632 
      WHEN  434 => wave := "001001111001"; --        633 
      WHEN  435 => wave := "001001111010"; --        634 
      WHEN  436 => wave := "001001111100"; --        636 
      WHEN  437 => wave := "001001111101"; --        637 
      WHEN  438 => wave := "001001111110"; --        638 
      WHEN  439 => wave := "001001111111"; --        639 
      WHEN  440 => wave := "001010000000"; --        640 
      WHEN  441 => wave := "001010000010"; --        642 
      WHEN  442 => wave := "001010000011"; --        643 
      WHEN  443 => wave := "001010000100"; --        644 
      WHEN  444 => wave := "001010000101"; --        645 
      WHEN  445 => wave := "001010000111"; --        647 
      WHEN  446 => wave := "001010001000"; --        648 
      WHEN  447 => wave := "001010001001"; --        649 
      WHEN  448 => wave := "001010001010"; --        650 
      WHEN  449 => wave := "001010001011"; --        651 
      WHEN  450 => wave := "001010001101"; --        653 
      WHEN  451 => wave := "001010001110"; --        654 
      WHEN  452 => wave := "001010001111"; --        655 
      WHEN  453 => wave := "001010010000"; --        656 
      WHEN  454 => wave := "001010010001"; --        657 
      WHEN  455 => wave := "001010010011"; --        659 
      WHEN  456 => wave := "001010010100"; --        660 
      WHEN  457 => wave := "001010010101"; --        661 
      WHEN  458 => wave := "001010010110"; --        662 
      WHEN  459 => wave := "001010010111"; --        663 
      WHEN  460 => wave := "001010011001"; --        665 
      WHEN  461 => wave := "001010011010"; --        666 
      WHEN  462 => wave := "001010011011"; --        667 
      WHEN  463 => wave := "001010011100"; --        668 
      WHEN  464 => wave := "001010011101"; --        669 
      WHEN  465 => wave := "001010011111"; --        671 
      WHEN  466 => wave := "001010100000"; --        672 
      WHEN  467 => wave := "001010100001"; --        673 
      WHEN  468 => wave := "001010100010"; --        674 
      WHEN  469 => wave := "001010100011"; --        675 
      WHEN  470 => wave := "001010100101"; --        677 
      WHEN  471 => wave := "001010100110"; --        678 
      WHEN  472 => wave := "001010100111"; --        679 
      WHEN  473 => wave := "001010101000"; --        680 
      WHEN  474 => wave := "001010101001"; --        681 
      WHEN  475 => wave := "001010101010"; --        682 
      WHEN  476 => wave := "001010101100"; --        684 
      WHEN  477 => wave := "001010101101"; --        685 
      WHEN  478 => wave := "001010101110"; --        686 
      WHEN  479 => wave := "001010101111"; --        687 
      WHEN  480 => wave := "001010110000"; --        688 
      WHEN  481 => wave := "001010110001"; --        689 
      WHEN  482 => wave := "001010110011"; --        691 
      WHEN  483 => wave := "001010110100"; --        692 
      WHEN  484 => wave := "001010110101"; --        693 
      WHEN  485 => wave := "001010110110"; --        694 
      WHEN  486 => wave := "001010110111"; --        695 
      WHEN  487 => wave := "001010111000"; --        696 
      WHEN  488 => wave := "001010111010"; --        698 
      WHEN  489 => wave := "001010111011"; --        699 
      WHEN  490 => wave := "001010111100"; --        700 
      WHEN  491 => wave := "001010111101"; --        701 
      WHEN  492 => wave := "001010111110"; --        702 
      WHEN  493 => wave := "001010111111"; --        703 
      WHEN  494 => wave := "001011000000"; --        704 
      WHEN  495 => wave := "001011000010"; --        706 
      WHEN  496 => wave := "001011000011"; --        707 
      WHEN  497 => wave := "001011000100"; --        708 
      WHEN  498 => wave := "001011000101"; --        709 
      WHEN  499 => wave := "001011000110"; --        710 
      WHEN  500 => wave := "001011000111"; --        711 
      WHEN  501 => wave := "001011001000"; --        712 
      WHEN  502 => wave := "001011001001"; --        713 
      WHEN  503 => wave := "001011001011"; --        715 
      WHEN  504 => wave := "001011001100"; --        716 
      WHEN  505 => wave := "001011001101"; --        717 
      WHEN  506 => wave := "001011001110"; --        718 
      WHEN  507 => wave := "001011001111"; --        719 
      WHEN  508 => wave := "001011010000"; --        720 
      WHEN  509 => wave := "001011010001"; --        721 
      WHEN  510 => wave := "001011010010"; --        722 
      WHEN OTHERS => wave := "001011010100"; --        724 
    END CASE; 

    sine <= wave; 

  END PROCESS; 
END ARCHITECTURE rtl; 
