LIBRARY IEEE; 
  USE IEEE.std_logic_1164.all; 
  USE IEEE.numeric_std.all; 

ENTITY COREFFT_C0_COREFFT_C0_0_twiddle IS 
  PORT ( 
    A : IN std_logic_vector(9 DOWNTO 0); 
    T : OUT std_logic_vector(47 DOWNTO 0)); 
END ENTITY COREFFT_C0_COREFFT_C0_0_twiddle; 

ARCHITECTURE rtl OF COREFFT_C0_COREFFT_C0_0_twiddle IS 
  SIGNAL A_int : integer; 
BEGIN 
  A_int <= to_integer(unsigned(A)); 
  PROCESS (A_int) 
    VARIABLE Ti  : std_logic_vector(47 DOWNTO 0); 
  BEGIN 
    CASE A_int IS      -- synopsys parallel_case     
      WHEN    0 => Ti := "000000000000000000000000011111111111111111111111"; --         +0   +8388607
      WHEN    1 => Ti := "111111111001101101111000011111111111111111011000"; --     -25736   +8388568
      WHEN    2 => Ti := "111111110011011011110000011111111111111101100001"; --     -51472   +8388449
      WHEN    3 => Ti := "111111101101001001101001011111111111111010011100"; --     -77207   +8388252
      WHEN    4 => Ti := "111111100110110111100011011111111111110110000111"; --    -102941   +8387975
      WHEN    5 => Ti := "111111100000100101011101011111111111110000100100"; --    -128675   +8387620
      WHEN    6 => Ti := "111111011010010011011001011111111111101001110010"; --    -154407   +8387186
      WHEN    7 => Ti := "111111010100000001010110011111111111100001110001"; --    -180138   +8386673
      WHEN    8 => Ti := "111111001101101111010101011111111111011000100001"; --    -205867   +8386081
      WHEN    9 => Ti := "111111000111011101010110011111111111001110000001"; --    -231594   +8385409
      WHEN   10 => Ti := "111111000001001011011001011111111111000010010011"; --    -257319   +8384659
      WHEN   11 => Ti := "111110111010111001011111011111111110110101010111"; --    -283041   +8383831
      WHEN   12 => Ti := "111110110100100111100111011111111110100111001011"; --    -308761   +8382923
      WHEN   13 => Ti := "111110101110010101110010011111111110010111110000"; --    -334478   +8381936
      WHEN   14 => Ti := "111110101000000100000000011111111110000111000110"; --    -360192   +8380870
      WHEN   15 => Ti := "111110100001110010010001011111111101110101001110"; --    -385903   +8379726
      WHEN   16 => Ti := "111110011011100000100111011111111101100010000111"; --    -411609   +8378503
      WHEN   17 => Ti := "111110010101001111000000011111111101001101110000"; --    -437312   +8377200
      WHEN   18 => Ti := "111110001110111101011101011111111100111000001011"; --    -463011   +8375819
      WHEN   19 => Ti := "111110001000101011111110011111111100100001010111"; --    -488706   +8374359
      WHEN   20 => Ti := "111110000010011010100100011111111100001001010101"; --    -514396   +8372821
      WHEN   21 => Ti := "111101111100001001001111011111111011110000000011"; --    -540081   +8371203
      WHEN   22 => Ti := "111101110101110111111111011111111011010101100011"; --    -565761   +8369507
      WHEN   23 => Ti := "111101101111100110110101011111111010111001110100"; --    -591435   +8367732
      WHEN   24 => Ti := "111101101001010101110000011111111010011100110110"; --    -617104   +8365878
      WHEN   25 => Ti := "111101100011000100110001011111111001111110101001"; --    -642767   +8363945
      WHEN   26 => Ti := "111101011100110011110111011111111001011111001110"; --    -668425   +8361934
      WHEN   27 => Ti := "111101010110100011000100011111111000111110100100"; --    -694076   +8359844
      WHEN   28 => Ti := "111101010000010010011000011111111000011100101011"; --    -719720   +8357675
      WHEN   29 => Ti := "111101001010000001110010011111110111111001100100"; --    -745358   +8355428
      WHEN   30 => Ti := "111101000011110001010100011111110111010101001110"; --    -770988   +8353102
      WHEN   31 => Ti := "111100111101100000111101011111110110101111101001"; --    -796611   +8350697
      WHEN   32 => Ti := "111100110111010000101101011111110110001000110110"; --    -822227   +8348214
      WHEN   33 => Ti := "111100110001000000100101011111110101100000110100"; --    -847835   +8345652
      WHEN   34 => Ti := "111100101010110000100101011111110100110111100011"; --    -873435   +8343011
      WHEN   35 => Ti := "111100100100100000101101011111110100001101000100"; --    -899027   +8340292
      WHEN   36 => Ti := "111100011110010000111101011111110011100001010111"; --    -924611   +8337495
      WHEN   37 => Ti := "111100011000000001010110011111110010110100011011"; --    -950186   +8334619
      WHEN   38 => Ti := "111100010001110001111001011111110010000110010001"; --    -975751   +8331665
      WHEN   39 => Ti := "111100001011100010100100011111110001010110111000"; --   -1001308   +8328632
      WHEN   40 => Ti := "111100000101010011011001011111110000100110010001"; --   -1026855   +8325521
      WHEN   41 => Ti := "111011111111000100010111011111101111110100011011"; --   -1052393   +8322331
      WHEN   42 => Ti := "111011111000110101100000011111101111000001010111"; --   -1077920   +8319063
      WHEN   43 => Ti := "111011110010100110110010011111101110001101000101"; --   -1103438   +8315717
      WHEN   44 => Ti := "111011101100011000001111011111101101010111100101"; --   -1128945   +8312293
      WHEN   45 => Ti := "111011100110001001110111011111101100100000110110"; --   -1154441   +8308790
      WHEN   46 => Ti := "111011011111111011101001011111101011101000111001"; --   -1179927   +8305209
      WHEN   47 => Ti := "111011011001101101100111011111101010101111101110"; --   -1205401   +8301550
      WHEN   48 => Ti := "111011010011011111110000011111101001110101010101"; --   -1230864   +8297813
      WHEN   49 => Ti := "111011001101010010000100011111101000111001101110"; --   -1256316   +8293998
      WHEN   50 => Ti := "111011000111000100100100011111100111111100111000"; --   -1281756   +8290104
      WHEN   51 => Ti := "111011000000110111010001011111100110111110110101"; --   -1307183   +8286133
      WHEN   52 => Ti := "111010111010101010001001011111100101111111100100"; --   -1332599   +8282084
      WHEN   53 => Ti := "111010110100011101001111011111100100111111000100"; --   -1358001   +8277956
      WHEN   54 => Ti := "111010101110010000100001011111100011111101010111"; --   -1383391   +8273751
      WHEN   55 => Ti := "111010101000000100000000011111100010111010011100"; --   -1408768   +8269468
      WHEN   56 => Ti := "111010100001110111101100011111100001110110010011"; --   -1434132   +8265107
      WHEN   57 => Ti := "111010011011101011100110011111100000110000111100"; --   -1459482   +8260668
      WHEN   58 => Ti := "111010010101011111101101011111011111101010011000"; --   -1484819   +8256152
      WHEN   59 => Ti := "111010001111010100000011011111011110100010100101"; --   -1510141   +8251557
      WHEN   60 => Ti := "111010001001001000100110011111011101011001100110"; --   -1535450   +8246886
      WHEN   61 => Ti := "111010000010111101011000011111011100001111011000"; --   -1560744   +8242136
      WHEN   62 => Ti := "111001111100110010011001011111011011000011111101"; --   -1586023   +8237309
      WHEN   63 => Ti := "111001110110100111101001011111011001110111010100"; --   -1611287   +8232404
      WHEN   64 => Ti := "111001110000011101001000011111011000101001011110"; --   -1636536   +8227422
      WHEN   65 => Ti := "111001101010010010110110011111010111011010011011"; --   -1661770   +8222363
      WHEN   66 => Ti := "111001100100001000110100011111010110001010001010"; --   -1686988   +8217226
      WHEN   67 => Ti := "111001011101111111000010011111010100111000101100"; --   -1712190   +8212012
      WHEN   68 => Ti := "111001010111110101100000011111010011100110000000"; --   -1737376   +8206720
      WHEN   69 => Ti := "111001010001101100001110011111010010010010000111"; --   -1762546   +8201351
      WHEN   70 => Ti := "111001001011100011001101011111010000111101000001"; --   -1787699   +8195905
      WHEN   71 => Ti := "111001000101011010011101011111001111100110101110"; --   -1812835   +8190382
      WHEN   72 => Ti := "111000111111010001111110011111001110001111001110"; --   -1837954   +8184782
      WHEN   73 => Ti := "111000111001001001110000011111001100110110100000"; --   -1863056   +8179104
      WHEN   74 => Ti := "111000110011000001110100011111001011011100100110"; --   -1888140   +8173350
      WHEN   75 => Ti := "111000101100111010001001011111001010000001011111"; --   -1913207   +8167519
      WHEN   76 => Ti := "111000100110110010110000011111001000100101001011"; --   -1938256   +8161611
      WHEN   77 => Ti := "111000100000101011101010011111000111000111101010"; --   -1963286   +8155626
      WHEN   78 => Ti := "111000011010100100110110011111000101101000111100"; --   -1988298   +8149564
      WHEN   79 => Ti := "111000010100011110010101011111000100001001000010"; --   -2013291   +8143426
      WHEN   80 => Ti := "111000001110011000000111011111000010100111111011"; --   -2038265   +8137211
      WHEN   81 => Ti := "111000001000010010001100011111000001000101100111"; --   -2063220   +8130919
      WHEN   82 => Ti := "111000000010001100100100011110111111100010000111"; --   -2088156   +8124551
      WHEN   83 => Ti := "110111111100000111010000011110111101111101011011"; --   -2113072   +8118107
      WHEN   84 => Ti := "110111110110000010010000011110111100010111100010"; --   -2137968   +8111586
      WHEN   85 => Ti := "110111101111111101100100011110111010110000011100"; --   -2162844   +8104988
      WHEN   86 => Ti := "110111101001111001001101011110111001001000001011"; --   -2187699   +8098315
      WHEN   87 => Ti := "110111100011110101001010011110110111011110101101"; --   -2212534   +8091565
      WHEN   88 => Ti := "110111011101110001011011011110110101110100000011"; --   -2237349   +8084739
      WHEN   89 => Ti := "110111010111101110000010011110110100001000001101"; --   -2262142   +8077837
      WHEN   90 => Ti := "110111010001101010111111011110110010011011001010"; --   -2286913   +8070858
      WHEN   91 => Ti := "110111001011101000010000011110110000101100111100"; --   -2311664   +8063804
      WHEN   92 => Ti := "110111000101100101111000011110101110111101100010"; --   -2336392   +8056674
      WHEN   93 => Ti := "110110111111100011110101011110101101001100111100"; --   -2361099   +8049468
      WHEN   94 => Ti := "110110111001100010001001011110101011011011001011"; --   -2385783   +8042187
      WHEN   95 => Ti := "110110110011100000110011011110101001101000001101"; --   -2410445   +8034829
      WHEN   96 => Ti := "110110101101011111110100011110100111110100000100"; --   -2435084   +8027396
      WHEN   97 => Ti := "110110100111011111001100011110100101111110110000"; --   -2459700   +8019888
      WHEN   98 => Ti := "110110100001011110111011011110100100001000010000"; --   -2484293   +8012304
      WHEN   99 => Ti := "110110011011011111000001011110100010010000100100"; --   -2508863   +8004644
      WHEN  100 => Ti := "110110010101011111011111011110100000010111101110"; --   -2533409   +7996910
      WHEN  101 => Ti := "110110001111100000010101011110011110011101101100"; --   -2557931   +7989100
      WHEN  102 => Ti := "110110001001100001100010011110011100100010011110"; --   -2582430   +7981214
      WHEN  103 => Ti := "110110000011100011001000011110011010100110000110"; --   -2606904   +7973254
      WHEN  104 => Ti := "110101111101100101000111011110011000101000100011"; --   -2631353   +7965219
      WHEN  105 => Ti := "110101110111100111011111011110010110101001110100"; --   -2655777   +7957108
      WHEN  106 => Ti := "110101110001101010001111011110010100101001111011"; --   -2680177   +7948923
      WHEN  107 => Ti := "110101101011101101011001011110010010101000110111"; --   -2704551   +7940663
      WHEN  108 => Ti := "110101100101110000111100011110010000100110101000"; --   -2728900   +7932328
      WHEN  109 => Ti := "110101011111110100111001011110001110100011001111"; --   -2753223   +7923919
      WHEN  110 => Ti := "110101011001111001001111011110001100011110101011"; --   -2777521   +7915435
      WHEN  111 => Ti := "110101010011111110000000011110001010011000111100"; --   -2801792   +7906876
      WHEN  112 => Ti := "110101001110000011001011011110001000010010000011"; --   -2826037   +7898243
      WHEN  113 => Ti := "110101001000001000110001011110000110001010000000"; --   -2850255   +7889536
      WHEN  114 => Ti := "110101000010001110110010011110000100000000110010"; --   -2874446   +7880754
      WHEN  115 => Ti := "110100111100010101001110011110000001110110011010"; --   -2898610   +7871898
      WHEN  116 => Ti := "110100110110011100000101011101111111101010111001"; --   -2922747   +7862969
      WHEN  117 => Ti := "110100110000100011010111011101111101011110001101"; --   -2946857   +7853965
      WHEN  118 => Ti := "110100101010101011000101011101111011010000010111"; --   -2970939   +7844887
      WHEN  119 => Ti := "110100100100110011010000011101111001000001010111"; --   -2994992   +7835735
      WHEN  120 => Ti := "110100011110111011110110011101110110110001001110"; --   -3019018   +7826510
      WHEN  121 => Ti := "110100011001000100111001011101110100011111111011"; --   -3043015   +7817211
      WHEN  122 => Ti := "110100010011001110011000011101110010001101011110"; --   -3066984   +7807838
      WHEN  123 => Ti := "110100001101011000010101011101101111111001111000"; --   -3090923   +7798392
      WHEN  124 => Ti := "110100000111100010101110011101101101100101001001"; --   -3114834   +7788873
      WHEN  125 => Ti := "110100000001101101100101011101101011001111010000"; --   -3138715   +7779280
      WHEN  126 => Ti := "110011111011111000111001011101101000111000001110"; --   -3162567   +7769614
      WHEN  127 => Ti := "110011110110000100101011011101100110100000000011"; --   -3186389   +7759875
      WHEN  128 => Ti := "110011110000010000111011011101100100000110101110"; --   -3210181   +7750062
      WHEN  129 => Ti := "110011101010011101101001011101100001101100010001"; --   -3233943   +7740177
      WHEN  130 => Ti := "110011100100101010110110011101011111010000101011"; --   -3257674   +7730219
      WHEN  131 => Ti := "110011011110111000100001011101011100110011111100"; --   -3281375   +7720188
      WHEN  132 => Ti := "110011011001000110101100011101011010010110000101"; --   -3305044   +7710085
      WHEN  133 => Ti := "110011010011010101010101011101010111110111000101"; --   -3328683   +7699909
      WHEN  134 => Ti := "110011001101100100011110011101010101010110111100"; --   -3352290   +7689660
      WHEN  135 => Ti := "110011000111110100000110011101010010110101101100"; --   -3375866   +7679340
      WHEN  136 => Ti := "110011000010000100001110011101010000010011010010"; --   -3399410   +7668946
      WHEN  137 => Ti := "110010111100010100110110011101001101101111110001"; --   -3422922   +7658481
      WHEN  138 => Ti := "110010110110100101111110011101001011001011001000"; --   -3446402   +7647944
      WHEN  139 => Ti := "110010110000110111100111011101001000100101010110"; --   -3469849   +7637334
      WHEN  140 => Ti := "110010101011001001110000011101000101111110011101"; --   -3493264   +7626653
      WHEN  141 => Ti := "110010100101011100011010011101000011010110011100"; --   -3516646   +7615900
      WHEN  142 => Ti := "110010011111101111100110011101000000101101010011"; --   -3539994   +7605075
      WHEN  143 => Ti := "110010011010000011010010011100111110000011000011"; --   -3563310   +7594179
      WHEN  144 => Ti := "110010010100010111100000011100111011010111101011"; --   -3586592   +7583211
      WHEN  145 => Ti := "110010001110101100010000011100111000101011001100"; --   -3609840   +7572172
      WHEN  146 => Ti := "110010001001000001100010011100110101111101100101"; --   -3633054   +7561061
      WHEN  147 => Ti := "110010000011010111010110011100110011001110111000"; --   -3656234   +7549880
      WHEN  148 => Ti := "110001111101101101101101011100110000011111000011"; --   -3679379   +7538627
      WHEN  149 => Ti := "110001111000000100100110011100101101101110000111"; --   -3702490   +7527303
      WHEN  150 => Ti := "110001110010011100000010011100101010111100000101"; --   -3725566   +7515909
      WHEN  151 => Ti := "110001101100110100000001011100101000001000111100"; --   -3748607   +7504444
      WHEN  152 => Ti := "110001100111001100100011011100100101010100101100"; --   -3771613   +7492908
      WHEN  153 => Ti := "110001100001100101101001011100100010011111010101"; --   -3794583   +7481301
      WHEN  154 => Ti := "110001011011111111010011011100011111101000111000"; --   -3817517   +7469624
      WHEN  155 => Ti := "110001010110011001100000011100011100110001010101"; --   -3840416   +7457877
      WHEN  156 => Ti := "110001010000110100010010011100011001111000101100"; --   -3863278   +7446060
      WHEN  157 => Ti := "110001001011001111101000011100010110111110111101"; --   -3886104   +7434173
      WHEN  158 => Ti := "110001000101101011100010011100010100000100000111"; --   -3908894   +7422215
      WHEN  159 => Ti := "110001000000001000000010011100010001001000001100"; --   -3931646   +7410188
      WHEN  160 => Ti := "110000111010100101000110011100001110001011001011"; --   -3954362   +7398091
      WHEN  161 => Ti := "110000110101000010110000011100001011001101000100"; --   -3977040   +7385924
      WHEN  162 => Ti := "110000101111100000111111011100001000001101111000"; --   -3999681   +7373688
      WHEN  163 => Ti := "110000101001111111110011011100000101001101100111"; --   -4022285   +7361383
      WHEN  164 => Ti := "110000100100011111001110011100000010001100010000"; --   -4044850   +7349008
      WHEN  165 => Ti := "110000011110111111001110011011111111001001110100"; --   -4067378   +7336564
      WHEN  166 => Ti := "110000011001011111110101011011111100000110010011"; --   -4089867   +7324051
      WHEN  167 => Ti := "110000010100000001000011011011111001000001101101"; --   -4112317   +7311469
      WHEN  168 => Ti := "110000001110100010110111011011110101111100000010"; --   -4134729   +7298818
      WHEN  169 => Ti := "110000001001000101010010011011110010110101010010"; --   -4157102   +7286098
      WHEN  170 => Ti := "110000000011101000010100011011101111101101011110"; --   -4179436   +7273310
      WHEN  171 => Ti := "101111111110001011111101011011101100100100100110"; --   -4201731   +7260454
      WHEN  172 => Ti := "101111111000110000001110011011101001011010101001"; --   -4223986   +7247529
      WHEN  173 => Ti := "101111110011010101000111011011100110001111101000"; --   -4246201   +7234536
      WHEN  174 => Ti := "101111101101111010101000011011100011000011100010"; --   -4268376   +7221474
      WHEN  175 => Ti := "101111101000100000110001011011011111110110011001"; --   -4290511   +7208345
      WHEN  176 => Ti := "101111100011000111100010011011011100101000001100"; --   -4312606   +7195148
      WHEN  177 => Ti := "101111011101101110111100011011011001011000111011"; --   -4334660   +7181883
      WHEN  178 => Ti := "101111011000010110111111011011010110001000100111"; --   -4356673   +7168551
      WHEN  179 => Ti := "101111010010111111101010011011010010110111001111"; --   -4378646   +7155151
      WHEN  180 => Ti := "101111001101101000111111011011001111100100110100"; --   -4400577   +7141684
      WHEN  181 => Ti := "101111001000010010111110011011001100010001010110"; --   -4422466   +7128150
      WHEN  182 => Ti := "101111000010111101100110011011001000111100110100"; --   -4444314   +7114548
      WHEN  183 => Ti := "101110111101101000110111011011000101100111010000"; --   -4466121   +7100880
      WHEN  184 => Ti := "101110111000010100110011011011000010010000101001"; --   -4487885   +7087145
      WHEN  185 => Ti := "101110110011000001011001011010111110111000111111"; --   -4509607   +7073343
      WHEN  186 => Ti := "101110101101101110101010011010111011100000010010"; --   -4531286   +7059474
      WHEN  187 => Ti := "101110101000011100100101011010111000000110100011"; --   -4552923   +7045539
      WHEN  188 => Ti := "101110100011001011001011011010110100101011110010"; --   -4574517   +7031538
      WHEN  189 => Ti := "101110011101111010011100011010110001001111111110"; --   -4596068   +7017470
      WHEN  190 => Ti := "101110011000101010011000011010101101110011001001"; --   -4617576   +7003337
      WHEN  191 => Ti := "101110010011011011000000011010101010010101010001"; --   -4639040   +6989137
      WHEN  192 => Ti := "101110001110001100010100011010100110110110011000"; --   -4660460   +6974872
      WHEN  193 => Ti := "101110001000111110010011011010100011010110011101"; --   -4681837   +6960541
      WHEN  194 => Ti := "101110000011110000111110011010011111110101100000"; --   -4703170   +6946144
      WHEN  195 => Ti := "101101111110100100010110011010011100010011100011"; --   -4724458   +6931683
      WHEN  196 => Ti := "101101111001011000011010011010011000110000100100"; --   -4745702   +6917156
      WHEN  197 => Ti := "101101110100001101001011011010010101001100100011"; --   -4766901   +6902563
      WHEN  198 => Ti := "101101101111000010101001011010010001100111100010"; --   -4788055   +6887906
      WHEN  199 => Ti := "101101101001111000110011011010001110000001100000"; --   -4809165   +6873184
      WHEN  200 => Ti := "101101100100101111101011011010001010011010011110"; --   -4830229   +6858398
      WHEN  201 => Ti := "101101011111100111010001011010000110110010011010"; --   -4851247   +6843546
      WHEN  202 => Ti := "101101011010011111100100011010000011001001010111"; --   -4872220   +6828631
      WHEN  203 => Ti := "101101010101011000100101011001111111011111010011"; --   -4893147   +6813651
      WHEN  204 => Ti := "101101010000010010010100011001111011110100001111"; --   -4914028   +6798607
      WHEN  205 => Ti := "101101001011001100110001011001111000001000001011"; --   -4934863   +6783499
      WHEN  206 => Ti := "101101000110000111111101011001110100011011000111"; --   -4955651   +6768327
      WHEN  207 => Ti := "101101000001000011110111011001110000101101000011"; --   -4976393   +6753091
      WHEN  208 => Ti := "101100111100000000100001011001101100111110000000"; --   -4997087   +6737792
      WHEN  209 => Ti := "101100110110111101111001011001101001001101111110"; --   -5017735   +6722430
      WHEN  210 => Ti := "101100110001111100000000011001100101011100111100"; --   -5038336   +6707004
      WHEN  211 => Ti := "101100101100111010110111011001100001101010111011"; --   -5058889   +6691515
      WHEN  212 => Ti := "101100100111111010011110011001011101110111111011"; --   -5079394   +6675963
      WHEN  213 => Ti := "101100100010111010110100011001011010000011111100"; --   -5099852   +6660348
      WHEN  214 => Ti := "101100011101111011111011011001010110001110111111"; --   -5120261   +6644671
      WHEN  215 => Ti := "101100011000111101110001011001010010011001000011"; --   -5140623   +6628931
      WHEN  216 => Ti := "101100010100000000011000011001001110100010001000"; --   -5160936   +6613128
      WHEN  217 => Ti := "101100001111000011101111011001001010101010010000"; --   -5181201   +6597264
      WHEN  218 => Ti := "101100001010000111111000011001000110110001011001"; --   -5201416   +6581337
      WHEN  219 => Ti := "101100000101001100110001011001000010110111100100"; --   -5221583   +6565348
      WHEN  220 => Ti := "101100000000010010011011011000111110111100110010"; --   -5241701   +6549298
      WHEN  221 => Ti := "101011111011011000110111011000111011000001000010"; --   -5261769   +6533186
      WHEN  222 => Ti := "101011110110100000000100011000110111000100010100"; --   -5281788   +6517012
      WHEN  223 => Ti := "101011110001101000000011011000110011000110101001"; --   -5301757   +6500777
      WHEN  224 => Ti := "101011101100110000110100011000101111001000000001"; --   -5321676   +6484481
      WHEN  225 => Ti := "101011100111111010010111011000101011001000011100"; --   -5341545   +6468124
      WHEN  226 => Ti := "101011100011000100101100011000100111000111111010"; --   -5361364   +6451706
      WHEN  227 => Ti := "101011011110001111110100011000100011000110011011"; --   -5381132   +6435227
      WHEN  228 => Ti := "101011011001011011101110011000011111000011111111"; --   -5400850   +6418687
      WHEN  229 => Ti := "101011010100101000011011011000011011000000101000"; --   -5420517   +6402088
      WHEN  230 => Ti := "101011001111110101111100011000010110111100010100"; --   -5440132   +6385428
      WHEN  231 => Ti := "101011001011000100001111011000010010110111000100"; --   -5459697   +6368708
      WHEN  232 => Ti := "101011000110010011010110011000001110110000110111"; --   -5479210   +6351927
      WHEN  233 => Ti := "101011000001100011010000011000001010101001110000"; --   -5498672   +6335088
      WHEN  234 => Ti := "101010111100110011111110011000000110100001101100"; --   -5518082   +6318188
      WHEN  235 => Ti := "101010111000000101100000011000000010011000101101"; --   -5537440   +6301229
      WHEN  236 => Ti := "101010110011010111110110010111111110001110110011"; --   -5556746   +6284211
      WHEN  237 => Ti := "101010101110101011000001010111111010000011111101"; --   -5575999   +6267133
      WHEN  238 => Ti := "101010101001111111000000010111110101111000001101"; --   -5595200   +6249997
      WHEN  239 => Ti := "101010100101010011110011010111110001101011100010"; --   -5614349   +6232802
      WHEN  240 => Ti := "101010100000101001011100010111101101011101111100"; --   -5633444   +6215548
      WHEN  241 => Ti := "101010011011111111111001010111101001001111011011"; --   -5652487   +6198235
      WHEN  242 => Ti := "101010010111010111001100010111100101000000000001"; --   -5671476   +6180865
      WHEN  243 => Ti := "101010010010101111010100010111100000101111101100"; --   -5690412   +6163436
      WHEN  244 => Ti := "101010001110001000010010010111011100011110011101"; --   -5709294   +6145949
      WHEN  245 => Ti := "101010001001100010000101010111011000001100010100"; --   -5728123   +6128404
      WHEN  246 => Ti := "101010000100111100101110010111010011111001010001"; --   -5746898   +6110801
      WHEN  247 => Ti := "101010000000011000001110010111001111100101010101"; --   -5765618   +6093141
      WHEN  248 => Ti := "101001111011110100100011010111001011010000100000"; --   -5784285   +6075424
      WHEN  249 => Ti := "101001110111010001101111010111000110111010110010"; --   -5802897   +6057650
      WHEN  250 => Ti := "101001110010101111110010010111000010100100001010"; --   -5821454   +6039818
      WHEN  251 => Ti := "101001101110001110101100010110111110001100101010"; --   -5839956   +6021930
      WHEN  252 => Ti := "101001101001101110011100010110111001110100010001"; --   -5858404   +6003985
      WHEN  253 => Ti := "101001100101001111000100010110110101011010111111"; --   -5876796   +5985983
      WHEN  254 => Ti := "101001100000110000100011010110110001000000110101"; --   -5895133   +5967925
      WHEN  255 => Ti := "101001011100010010111001010110101100100101110011"; --   -5913415   +5949811
      WHEN  256 => Ti := "101001010111110110000111010110101000001001111001"; --   -5931641   +5931641
      WHEN  257 => Ti := "101001010011011010001101010110100011101101000111"; --   -5949811   +5913415
      WHEN  258 => Ti := "101001001110111111001011010110011111001111011101"; --   -5967925   +5895133
      WHEN  259 => Ti := "101001001010100101000001010110011010110000111100"; --   -5985983   +5876796
      WHEN  260 => Ti := "101001000110001011101111010110010110010001100100"; --   -6003985   +5858404
      WHEN  261 => Ti := "101001000001110011010110010110010001110001010100"; --   -6021930   +5839956
      WHEN  262 => Ti := "101000111101011011110110010110001101010000001110"; --   -6039818   +5821454
      WHEN  263 => Ti := "101000111001000101001110010110001000101110010001"; --   -6057650   +5802897
      WHEN  264 => Ti := "101000110100101111100000010110000100001011011101"; --   -6075424   +5784285
      WHEN  265 => Ti := "101000110000011010101011010101111111100111110010"; --   -6093141   +5765618
      WHEN  266 => Ti := "101000101100000110101111010101111011000011010010"; --   -6110801   +5746898
      WHEN  267 => Ti := "101000100111110011101100010101110110011101111011"; --   -6128404   +5728123
      WHEN  268 => Ti := "101000100011100001100011010101110001110111101110"; --   -6145949   +5709294
      WHEN  269 => Ti := "101000011111010000010100010101101101010000101100"; --   -6163436   +5690412
      WHEN  270 => Ti := "101000011010111111111111010101101000101000110100"; --   -6180865   +5671476
      WHEN  271 => Ti := "101000010110110000100101010101100100000000000111"; --   -6198235   +5652487
      WHEN  272 => Ti := "101000010010100010000100010101011111010110100100"; --   -6215548   +5633444
      WHEN  273 => Ti := "101000001110010100011110010101011010101100001101"; --   -6232802   +5614349
      WHEN  274 => Ti := "101000001010000111110011010101010110000001000000"; --   -6249997   +5595200
      WHEN  275 => Ti := "101000000101111100000011010101010001010100111111"; --   -6267133   +5575999
      WHEN  276 => Ti := "101000000001110001001101010101001100101000001010"; --   -6284211   +5556746
      WHEN  277 => Ti := "100111111101100111010011010101000111111010100000"; --   -6301229   +5537440
      WHEN  278 => Ti := "100111111001011110010100010101000011001100000010"; --   -6318188   +5518082
      WHEN  279 => Ti := "100111110101010110010000010100111110011100110000"; --   -6335088   +5498672
      WHEN  280 => Ti := "100111110001001111001001010100111001101100101010"; --   -6351927   +5479210
      WHEN  281 => Ti := "100111101101001000111100010100110100111011110001"; --   -6368708   +5459697
      WHEN  282 => Ti := "100111101001000011101100010100110000001010000100"; --   -6385428   +5440132
      WHEN  283 => Ti := "100111100100111111011000010100101011010111100101"; --   -6402088   +5420517
      WHEN  284 => Ti := "100111100000111100000001010100100110100100010010"; --   -6418687   +5400850
      WHEN  285 => Ti := "100111011100111001100101010100100001110000001100"; --   -6435227   +5381132
      WHEN  286 => Ti := "100111011000111000000110010100011100111011010100"; --   -6451706   +5361364
      WHEN  287 => Ti := "100111010100110111100100010100011000000101101001"; --   -6468124   +5341545
      WHEN  288 => Ti := "100111010000110111111111010100010011001111001100"; --   -6484481   +5321676
      WHEN  289 => Ti := "100111001100111001010111010100001110010111111101"; --   -6500777   +5301757
      WHEN  290 => Ti := "100111001000111011101100010100001001011111111100"; --   -6517012   +5281788
      WHEN  291 => Ti := "100111000100111110111110010100000100100111001001"; --   -6533186   +5261769
      WHEN  292 => Ti := "100111000001000011001110010011111111101101100101"; --   -6549298   +5241701
      WHEN  293 => Ti := "100110111101001000011100010011111010110011001111"; --   -6565348   +5221583
      WHEN  294 => Ti := "100110111001001110100111010011110101111000001000"; --   -6581337   +5201416
      WHEN  295 => Ti := "100110110101010101110000010011110000111100010001"; --   -6597264   +5181201
      WHEN  296 => Ti := "100110110001011101111000010011101011111111101000"; --   -6613128   +5160936
      WHEN  297 => Ti := "100110101101100110111101010011100111000010001111"; --   -6628931   +5140623
      WHEN  298 => Ti := "100110101001110001000001010011100010000100000101"; --   -6644671   +5120261
      WHEN  299 => Ti := "100110100101111100000100010011011101000101001100"; --   -6660348   +5099852
      WHEN  300 => Ti := "100110100010001000000101010011011000000101100010"; --   -6675963   +5079394
      WHEN  301 => Ti := "100110011110010101000101010011010011000101001001"; --   -6691515   +5058889
      WHEN  302 => Ti := "100110011010100011000100010011001110000100000000"; --   -6707004   +5038336
      WHEN  303 => Ti := "100110010110110010000010010011001001000010000111"; --   -6722430   +5017735
      WHEN  304 => Ti := "100110010011000010000000010011000011111111011111"; --   -6737792   +4997087
      WHEN  305 => Ti := "100110001111010010111101010010111110111100001001"; --   -6753091   +4976393
      WHEN  306 => Ti := "100110001011100100111001010010111001111000000011"; --   -6768327   +4955651
      WHEN  307 => Ti := "100110000111110111110101010010110100110011001111"; --   -6783499   +4934863
      WHEN  308 => Ti := "100110000100001011110001010010101111101101101100"; --   -6798607   +4914028
      WHEN  309 => Ti := "100110000000100000101101010010101010100111011011"; --   -6813651   +4893147
      WHEN  310 => Ti := "100101111100110110101001010010100101100000011100"; --   -6828631   +4872220
      WHEN  311 => Ti := "100101111001001101100110010010100000011000101111"; --   -6843546   +4851247
      WHEN  312 => Ti := "100101110101100101100010010010011011010000010101"; --   -6858398   +4830229
      WHEN  313 => Ti := "100101110001111110100000010010010110000111001101"; --   -6873184   +4809165
      WHEN  314 => Ti := "100101101110011000011110010010010000111101010111"; --   -6887906   +4788055
      WHEN  315 => Ti := "100101101010110011011101010010001011110010110101"; --   -6902563   +4766901
      WHEN  316 => Ti := "100101100111001111011100010010000110100111100110"; --   -6917156   +4745702
      WHEN  317 => Ti := "100101100011101100011101010010000001011011101010"; --   -6931683   +4724458
      WHEN  318 => Ti := "100101100000001010100000010001111100001111000010"; --   -6946144   +4703170
      WHEN  319 => Ti := "100101011100101001100011010001110111000001101101"; --   -6960541   +4681837
      WHEN  320 => Ti := "100101011001001001101000010001110001110011101100"; --   -6974872   +4660460
      WHEN  321 => Ti := "100101010101101010101111010001101100100101000000"; --   -6989137   +4639040
      WHEN  322 => Ti := "100101010010001100110111010001100111010101101000"; --   -7003337   +4617576
      WHEN  323 => Ti := "100101001110110000000010010001100010000101100100"; --   -7017470   +4596068
      WHEN  324 => Ti := "100101001011010100001110010001011100110100110101"; --   -7031538   +4574517
      WHEN  325 => Ti := "100101000111111001011101010001010111100011011011"; --   -7045539   +4552923
      WHEN  326 => Ti := "100101000100011111101110010001010010010001010110"; --   -7059474   +4531286
      WHEN  327 => Ti := "100101000001000111000001010001001100111110100111"; --   -7073343   +4509607
      WHEN  328 => Ti := "100100111101101111010111010001000111101011001101"; --   -7087145   +4487885
      WHEN  329 => Ti := "100100111010011000110000010001000010010111001001"; --   -7100880   +4466121
      WHEN  330 => Ti := "100100110111000011001100010000111101000010011010"; --   -7114548   +4444314
      WHEN  331 => Ti := "100100110011101110101010010000110111101101000010"; --   -7128150   +4422466
      WHEN  332 => Ti := "100100110000011011001100010000110010010111000001"; --   -7141684   +4400577
      WHEN  333 => Ti := "100100101101001000110001010000101101000000010110"; --   -7155151   +4378646
      WHEN  334 => Ti := "100100101001110111011001010000100111101001000001"; --   -7168551   +4356673
      WHEN  335 => Ti := "100100100110100111000101010000100010010001000100"; --   -7181883   +4334660
      WHEN  336 => Ti := "100100100011010111110100010000011100111000011110"; --   -7195148   +4312606
      WHEN  337 => Ti := "100100100000001001100111010000010111011111001111"; --   -7208345   +4290511
      WHEN  338 => Ti := "100100011100111100011110010000010010000101011000"; --   -7221474   +4268376
      WHEN  339 => Ti := "100100011001110000011000010000001100101010111001"; --   -7234536   +4246201
      WHEN  340 => Ti := "100100010110100101010111010000000111001111110010"; --   -7247529   +4223986
      WHEN  341 => Ti := "100100010011011011011010010000000001110100000011"; --   -7260454   +4201731
      WHEN  342 => Ti := "100100010000010010100010001111111100010111101100"; --   -7273310   +4179436
      WHEN  343 => Ti := "100100001101001010101110001111110110111010101110"; --   -7286098   +4157102
      WHEN  344 => Ti := "100100001010000011111110001111110001011101001001"; --   -7298818   +4134729
      WHEN  345 => Ti := "100100000110111110010011001111101011111110111101"; --   -7311469   +4112317
      WHEN  346 => Ti := "100100000011111001101101001111100110100000001011"; --   -7324051   +4089867
      WHEN  347 => Ti := "100100000000110110001100001111100001000000110010"; --   -7336564   +4067378
      WHEN  348 => Ti := "100011111101110011110000001111011011100000110010"; --   -7349008   +4044850
      WHEN  349 => Ti := "100011111010110010011001001111010110000000001101"; --   -7361383   +4022285
      WHEN  350 => Ti := "100011110111110010001000001111010000011111000001"; --   -7373688   +3999681
      WHEN  351 => Ti := "100011110100110010111100001111001010111101010000"; --   -7385924   +3977040
      WHEN  352 => Ti := "100011110001110100110101001111000101011010111010"; --   -7398091   +3954362
      WHEN  353 => Ti := "100011101110110111110100001110111111110111111110"; --   -7410188   +3931646
      WHEN  354 => Ti := "100011101011111011111001001110111010010100011110"; --   -7422215   +3908894
      WHEN  355 => Ti := "100011101001000001000011001110110100110000011000"; --   -7434173   +3886104
      WHEN  356 => Ti := "100011100110000111010100001110101111001011101110"; --   -7446060   +3863278
      WHEN  357 => Ti := "100011100011001110101011001110101001100110100000"; --   -7457877   +3840416
      WHEN  358 => Ti := "100011100000010111001000001110100100000000101101"; --   -7469624   +3817517
      WHEN  359 => Ti := "100011011101100000101011001110011110011010010111"; --   -7481301   +3794583
      WHEN  360 => Ti := "100011011010101011010100001110011000110011011101"; --   -7492908   +3771613
      WHEN  361 => Ti := "100011010111110111000100001110010011001011111111"; --   -7504444   +3748607
      WHEN  362 => Ti := "100011010101000011111011001110001101100011111110"; --   -7515909   +3725566
      WHEN  363 => Ti := "100011010010010001111001001110000111111011011010"; --   -7527303   +3702490
      WHEN  364 => Ti := "100011001111100000111101001110000010010010010011"; --   -7538627   +3679379
      WHEN  365 => Ti := "100011001100110001001000001101111100101000101010"; --   -7549880   +3656234
      WHEN  366 => Ti := "100011001010000010011011001101110110111110011110"; --   -7561061   +3633054
      WHEN  367 => Ti := "100011000111010100110100001101110001010011110000"; --   -7572172   +3609840
      WHEN  368 => Ti := "100011000100101000010101001101101011101000100000"; --   -7583211   +3586592
      WHEN  369 => Ti := "100011000001111100111101001101100101111100101110"; --   -7594179   +3563310
      WHEN  370 => Ti := "100010111111010010101101001101100000010000011010"; --   -7605075   +3539994
      WHEN  371 => Ti := "100010111100101001100100001101011010100011100110"; --   -7615900   +3516646
      WHEN  372 => Ti := "100010111010000001100011001101010100110110010000"; --   -7626653   +3493264
      WHEN  373 => Ti := "100010110111011010101010001101001111001000011001"; --   -7637334   +3469849
      WHEN  374 => Ti := "100010110100110100111000001101001001011010000010"; --   -7647944   +3446402
      WHEN  375 => Ti := "100010110010010000001111001101000011101011001010"; --   -7658481   +3422922
      WHEN  376 => Ti := "100010101111101100101110001100111101111011110010"; --   -7668946   +3399410
      WHEN  377 => Ti := "100010101101001010010100001100111000001011111010"; --   -7679340   +3375866
      WHEN  378 => Ti := "100010101010101001000100001100110010011011100010"; --   -7689660   +3352290
      WHEN  379 => Ti := "100010101000001000111011001100101100101010101011"; --   -7699909   +3328683
      WHEN  380 => Ti := "100010100101101001111011001100100110111001010100"; --   -7710085   +3305044
      WHEN  381 => Ti := "100010100011001100000100001100100001000111011111"; --   -7720188   +3281375
      WHEN  382 => Ti := "100010100000101111010101001100011011010101001010"; --   -7730219   +3257674
      WHEN  383 => Ti := "100010011110010011101111001100010101100010010111"; --   -7740177   +3233943
      WHEN  384 => Ti := "100010011011111001010010001100001111101111000101"; --   -7750062   +3210181
      WHEN  385 => Ti := "100010011001011111111101001100001001111011010101"; --   -7759875   +3186389
      WHEN  386 => Ti := "100010010111000111110010001100000100000111000111"; --   -7769614   +3162567
      WHEN  387 => Ti := "100010010100110000110000001011111110010010011011"; --   -7779280   +3138715
      WHEN  388 => Ti := "100010010010011010110111001011111000011101010010"; --   -7788873   +3114834
      WHEN  389 => Ti := "100010010000000110001000001011110010100111101011"; --   -7798392   +3090923
      WHEN  390 => Ti := "100010001101110010100010001011101100110001101000"; --   -7807838   +3066984
      WHEN  391 => Ti := "100010001011100000000101001011100110111011000111"; --   -7817211   +3043015
      WHEN  392 => Ti := "100010001001001110110010001011100001000100001010"; --   -7826510   +3019018
      WHEN  393 => Ti := "100010000110111110101001001011011011001100110000"; --   -7835735   +2994992
      WHEN  394 => Ti := "100010000100101111101001001011010101010100111011"; --   -7844887   +2970939
      WHEN  395 => Ti := "100010000010100001110011001011001111011100101001"; --   -7853965   +2946857
      WHEN  396 => Ti := "100010000000010101000111001011001001100011111011"; --   -7862969   +2922747
      WHEN  397 => Ti := "100001111110001001100110001011000011101010110010"; --   -7871898   +2898610
      WHEN  398 => Ti := "100001111011111111001110001010111101110001001110"; --   -7880754   +2874446
      WHEN  399 => Ti := "100001111001110110000000001010110111110111001111"; --   -7889536   +2850255
      WHEN  400 => Ti := "100001110111101101111101001010110001111100110101"; --   -7898243   +2826037
      WHEN  401 => Ti := "100001110101100111000100001010101100000010000000"; --   -7906876   +2801792
      WHEN  402 => Ti := "100001110011100001010101001010100110000110110001"; --   -7915435   +2777521
      WHEN  403 => Ti := "100001110001011100110001001010100000001011000111"; --   -7923919   +2753223
      WHEN  404 => Ti := "100001101111011001011000001010011010001111000100"; --   -7932328   +2728900
      WHEN  405 => Ti := "100001101101010111001001001010010100010010100111"; --   -7940663   +2704551
      WHEN  406 => Ti := "100001101011010110000101001010001110010101110001"; --   -7948923   +2680177
      WHEN  407 => Ti := "100001101001010110001100001010001000011000100001"; --   -7957108   +2655777
      WHEN  408 => Ti := "100001100111010111011101001010000010011010111001"; --   -7965219   +2631353
      WHEN  409 => Ti := "100001100101011001111010001001111100011100111000"; --   -7973254   +2606904
      WHEN  410 => Ti := "100001100011011101100010001001110110011110011110"; --   -7981214   +2582430
      WHEN  411 => Ti := "100001100001100010010100001001110000011111101011"; --   -7989100   +2557931
      WHEN  412 => Ti := "100001011111101000010010001001101010100000100001"; --   -7996910   +2533409
      WHEN  413 => Ti := "100001011101101111011100001001100100100000111111"; --   -8004644   +2508863
      WHEN  414 => Ti := "100001011011110111110000001001011110100001000101"; --   -8012304   +2484293
      WHEN  415 => Ti := "100001011010000001010000001001011000100000110100"; --   -8019888   +2459700
      WHEN  416 => Ti := "100001011000001011111100001001010010100000001100"; --   -8027396   +2435084
      WHEN  417 => Ti := "100001010110010111110011001001001100011111001101"; --   -8034829   +2410445
      WHEN  418 => Ti := "100001010100100100110101001001000110011101110111"; --   -8042187   +2385783
      WHEN  419 => Ti := "100001010010110011000100001001000000011100001011"; --   -8049468   +2361099
      WHEN  420 => Ti := "100001010001000010011110001000111010011010001000"; --   -8056674   +2336392
      WHEN  421 => Ti := "100001001111010011000100001000110100010111110000"; --   -8063804   +2311664
      WHEN  422 => Ti := "100001001101100100110110001000101110010101000001"; --   -8070858   +2286913
      WHEN  423 => Ti := "100001001011110111110011001000101000010001111110"; --   -8077837   +2262142
      WHEN  424 => Ti := "100001001010001011111101001000100010001110100101"; --   -8084739   +2237349
      WHEN  425 => Ti := "100001001000100001010011001000011100001010110110"; --   -8091565   +2212534
      WHEN  426 => Ti := "100001000110110111110101001000010110000110110011"; --   -8098315   +2187699
      WHEN  427 => Ti := "100001000101001111100100001000010000000010011100"; --   -8104988   +2162844
      WHEN  428 => Ti := "100001000011101000011110001000001001111101110000"; --   -8111586   +2137968
      WHEN  429 => Ti := "100001000010000010100101001000000011111000110000"; --   -8118107   +2113072
      WHEN  430 => Ti := "100001000000011101111001000111111101110011011100"; --   -8124551   +2088156
      WHEN  431 => Ti := "100000111110111010011001000111110111101101110100"; --   -8130919   +2063220
      WHEN  432 => Ti := "100000111101011000000101000111110001100111111001"; --   -8137211   +2038265
      WHEN  433 => Ti := "100000111011110110111110000111101011100001101011"; --   -8143426   +2013291
      WHEN  434 => Ti := "100000111010010111000100000111100101011011001010"; --   -8149564   +1988298
      WHEN  435 => Ti := "100000111000111000010110000111011111010100010110"; --   -8155626   +1963286
      WHEN  436 => Ti := "100000110111011010110101000111011001001101010000"; --   -8161611   +1938256
      WHEN  437 => Ti := "100000110101111110100001000111010011000101110111"; --   -8167519   +1913207
      WHEN  438 => Ti := "100000110100100011011010000111001100111110001100"; --   -8173350   +1888140
      WHEN  439 => Ti := "100000110011001001100000000111000110110110010000"; --   -8179104   +1863056
      WHEN  440 => Ti := "100000110001110000110010000111000000101110000010"; --   -8184782   +1837954
      WHEN  441 => Ti := "100000110000011001010010000110111010100101100011"; --   -8190382   +1812835
      WHEN  442 => Ti := "100000101111000010111111000110110100011100110011"; --   -8195905   +1787699
      WHEN  443 => Ti := "100000101101101101111001000110101110010011110010"; --   -8201351   +1762546
      WHEN  444 => Ti := "100000101100011010000000000110101000001010100000"; --   -8206720   +1737376
      WHEN  445 => Ti := "100000101011000111010100000110100010000000111110"; --   -8212012   +1712190
      WHEN  446 => Ti := "100000101001110101110110000110011011110111001100"; --   -8217226   +1686988
      WHEN  447 => Ti := "100000101000100101100101000110010101101101001010"; --   -8222363   +1661770
      WHEN  448 => Ti := "100000100111010110100010000110001111100010111000"; --   -8227422   +1636536
      WHEN  449 => Ti := "100000100110001000101100000110001001011000010111"; --   -8232404   +1611287
      WHEN  450 => Ti := "100000100100111100000011000110000011001101100111"; --   -8237309   +1586023
      WHEN  451 => Ti := "100000100011110000101000000101111101000010101000"; --   -8242136   +1560744
      WHEN  452 => Ti := "100000100010100110011010000101110110110111011010"; --   -8246886   +1535450
      WHEN  453 => Ti := "100000100001011101011011000101110000101011111101"; --   -8251557   +1510141
      WHEN  454 => Ti := "100000100000010101101000000101101010100000010011"; --   -8256152   +1484819
      WHEN  455 => Ti := "100000011111001111000100000101100100010100011010"; --   -8260668   +1459482
      WHEN  456 => Ti := "100000011110001001101101000101011110001000010100"; --   -8265107   +1434132
      WHEN  457 => Ti := "100000011101000101100100000101010111111100000000"; --   -8269468   +1408768
      WHEN  458 => Ti := "100000011100000010101001000101010001101111011111"; --   -8273751   +1383391
      WHEN  459 => Ti := "100000011011000000111100000101001011100010110001"; --   -8277956   +1358001
      WHEN  460 => Ti := "100000011010000000011100000101000101010101110111"; --   -8282084   +1332599
      WHEN  461 => Ti := "100000011001000001001011000100111111001000101111"; --   -8286133   +1307183
      WHEN  462 => Ti := "100000011000000011001000000100111000111011011100"; --   -8290104   +1281756
      WHEN  463 => Ti := "100000010111000110010010000100110010101101111100"; --   -8293998   +1256316
      WHEN  464 => Ti := "100000010110001010101011000100101100100000010000"; --   -8297813   +1230864
      WHEN  465 => Ti := "100000010101010000010010000100100110010010011001"; --   -8301550   +1205401
      WHEN  466 => Ti := "100000010100010111000111000100100000000100010111"; --   -8305209   +1179927
      WHEN  467 => Ti := "100000010011011111001010000100011001110110001001"; --   -8308790   +1154441
      WHEN  468 => Ti := "100000010010101000011011000100010011100111110001"; --   -8312293   +1128945
      WHEN  469 => Ti := "100000010001110010111011000100001101011001001110"; --   -8315717   +1103438
      WHEN  470 => Ti := "100000010000111110101001000100000111001010100000"; --   -8319063   +1077920
      WHEN  471 => Ti := "100000010000001011100101000100000000111011101001"; --   -8322331   +1052393
      WHEN  472 => Ti := "100000001111011001101111000011111010101100100111"; --   -8325521   +1026855
      WHEN  473 => Ti := "100000001110101001001000000011110100011101011100"; --   -8328632   +1001308
      WHEN  474 => Ti := "100000001101111001101111000011101110001110000111"; --   -8331665    +975751
      WHEN  475 => Ti := "100000001101001011100101000011100111111110101010"; --   -8334619    +950186
      WHEN  476 => Ti := "100000001100011110101001000011100001101111000011"; --   -8337495    +924611
      WHEN  477 => Ti := "100000001011110010111100000011011011011111010011"; --   -8340292    +899027
      WHEN  478 => Ti := "100000001011001000011101000011010101001111011011"; --   -8343011    +873435
      WHEN  479 => Ti := "100000001010011111001100000011001110111111011011"; --   -8345652    +847835
      WHEN  480 => Ti := "100000001001110111001010000011001000101111010011"; --   -8348214    +822227
      WHEN  481 => Ti := "100000001001010000010111000011000010011111000011"; --   -8350697    +796611
      WHEN  482 => Ti := "100000001000101010110010000010111100001110101100"; --   -8353102    +770988
      WHEN  483 => Ti := "100000001000000110011100000010110101111110001110"; --   -8355428    +745358
      WHEN  484 => Ti := "100000000111100011010101000010101111101101101000"; --   -8357675    +719720
      WHEN  485 => Ti := "100000000111000001011100000010101001011100111100"; --   -8359844    +694076
      WHEN  486 => Ti := "100000000110100000110010000010100011001100001001"; --   -8361934    +668425
      WHEN  487 => Ti := "100000000110000001010111000010011100111011001111"; --   -8363945    +642767
      WHEN  488 => Ti := "100000000101100011001010000010010110101010010000"; --   -8365878    +617104
      WHEN  489 => Ti := "100000000101000110001100000010010000011001001011"; --   -8367732    +591435
      WHEN  490 => Ti := "100000000100101010011101000010001010001000000001"; --   -8369507    +565761
      WHEN  491 => Ti := "100000000100001111111101000010000011110110110001"; --   -8371203    +540081
      WHEN  492 => Ti := "100000000011110110101011000001111101100101011100"; --   -8372821    +514396
      WHEN  493 => Ti := "100000000011011110101001000001110111010100000010"; --   -8374359    +488706
      WHEN  494 => Ti := "100000000011000111110101000001110001000010100011"; --   -8375819    +463011
      WHEN  495 => Ti := "100000000010110010010000000001101010110001000000"; --   -8377200    +437312
      WHEN  496 => Ti := "100000000010011101111001000001100100011111011001"; --   -8378503    +411609
      WHEN  497 => Ti := "100000000010001010110010000001011110001101101111"; --   -8379726    +385903
      WHEN  498 => Ti := "100000000001111000111010000001010111111100000000"; --   -8380870    +360192
      WHEN  499 => Ti := "100000000001101000010000000001010001101010001110"; --   -8381936    +334478
      WHEN  500 => Ti := "100000000001011000110101000001001011011000011001"; --   -8382923    +308761
      WHEN  501 => Ti := "100000000001001010101001000001000101000110100001"; --   -8383831    +283041
      WHEN  502 => Ti := "100000000000111101101101000000111110110100100111"; --   -8384659    +257319
      WHEN  503 => Ti := "100000000000110001111111000000111000100010101010"; --   -8385409    +231594
      WHEN  504 => Ti := "100000000000100111011111000000110010010000101011"; --   -8386081    +205867
      WHEN  505 => Ti := "100000000000011110001111000000101011111110101010"; --   -8386673    +180138
      WHEN  506 => Ti := "100000000000010110001110000000100101101100100111"; --   -8387186    +154407
      WHEN  507 => Ti := "100000000000001111011100000000011111011010100011"; --   -8387620    +128675
      WHEN  508 => Ti := "100000000000001001111001000000011001001000011101"; --   -8387975    +102941
      WHEN  509 => Ti := "100000000000000101100100000000010010110110010111"; --   -8388252     +77207
      WHEN  510 => Ti := "100000000000000010011111000000001100100100010000"; --   -8388449     +51472
      WHEN  511 => Ti := "100000000000000000101000000000000110010010001000"; --   -8388568     +25736
      WHEN  512 => Ti := "100000000000000000000001000000000000000000000000"; --   -8388607         +0
      WHEN  513 => Ti := "100000000000000000101000111111111001101101111000"; --   -8388568     -25736
      WHEN  514 => Ti := "100000000000000010011111111111110011011011110000"; --   -8388449     -51472
      WHEN  515 => Ti := "100000000000000101100100111111101101001001101001"; --   -8388252     -77207
      WHEN  516 => Ti := "100000000000001001111001111111100110110111100011"; --   -8387975    -102941
      WHEN  517 => Ti := "100000000000001111011100111111100000100101011101"; --   -8387620    -128675
      WHEN  518 => Ti := "100000000000010110001110111111011010010011011001"; --   -8387186    -154407
      WHEN  519 => Ti := "100000000000011110001111111111010100000001010110"; --   -8386673    -180138
      WHEN  520 => Ti := "100000000000100111011111111111001101101111010101"; --   -8386081    -205867
      WHEN  521 => Ti := "100000000000110001111111111111000111011101010110"; --   -8385409    -231594
      WHEN  522 => Ti := "100000000000111101101101111111000001001011011001"; --   -8384659    -257319
      WHEN  523 => Ti := "100000000001001010101001111110111010111001011111"; --   -8383831    -283041
      WHEN  524 => Ti := "100000000001011000110101111110110100100111100111"; --   -8382923    -308761
      WHEN  525 => Ti := "100000000001101000010000111110101110010101110010"; --   -8381936    -334478
      WHEN  526 => Ti := "100000000001111000111010111110101000000100000000"; --   -8380870    -360192
      WHEN  527 => Ti := "100000000010001010110010111110100001110010010001"; --   -8379726    -385903
      WHEN  528 => Ti := "100000000010011101111001111110011011100000100111"; --   -8378503    -411609
      WHEN  529 => Ti := "100000000010110010010000111110010101001111000000"; --   -8377200    -437312
      WHEN  530 => Ti := "100000000011000111110101111110001110111101011101"; --   -8375819    -463011
      WHEN  531 => Ti := "100000000011011110101001111110001000101011111110"; --   -8374359    -488706
      WHEN  532 => Ti := "100000000011110110101011111110000010011010100100"; --   -8372821    -514396
      WHEN  533 => Ti := "100000000100001111111101111101111100001001001111"; --   -8371203    -540081
      WHEN  534 => Ti := "100000000100101010011101111101110101110111111111"; --   -8369507    -565761
      WHEN  535 => Ti := "100000000101000110001100111101101111100110110101"; --   -8367732    -591435
      WHEN  536 => Ti := "100000000101100011001010111101101001010101110000"; --   -8365878    -617104
      WHEN  537 => Ti := "100000000110000001010111111101100011000100110001"; --   -8363945    -642767
      WHEN  538 => Ti := "100000000110100000110010111101011100110011110111"; --   -8361934    -668425
      WHEN  539 => Ti := "100000000111000001011100111101010110100011000100"; --   -8359844    -694076
      WHEN  540 => Ti := "100000000111100011010101111101010000010010011000"; --   -8357675    -719720
      WHEN  541 => Ti := "100000001000000110011100111101001010000001110010"; --   -8355428    -745358
      WHEN  542 => Ti := "100000001000101010110010111101000011110001010100"; --   -8353102    -770988
      WHEN  543 => Ti := "100000001001010000010111111100111101100000111101"; --   -8350697    -796611
      WHEN  544 => Ti := "100000001001110111001010111100110111010000101101"; --   -8348214    -822227
      WHEN  545 => Ti := "100000001010011111001100111100110001000000100101"; --   -8345652    -847835
      WHEN  546 => Ti := "100000001011001000011101111100101010110000100101"; --   -8343011    -873435
      WHEN  547 => Ti := "100000001011110010111100111100100100100000101101"; --   -8340292    -899027
      WHEN  548 => Ti := "100000001100011110101001111100011110010000111101"; --   -8337495    -924611
      WHEN  549 => Ti := "100000001101001011100101111100011000000001010110"; --   -8334619    -950186
      WHEN  550 => Ti := "100000001101111001101111111100010001110001111001"; --   -8331665    -975751
      WHEN  551 => Ti := "100000001110101001001000111100001011100010100100"; --   -8328632   -1001308
      WHEN  552 => Ti := "100000001111011001101111111100000101010011011001"; --   -8325521   -1026855
      WHEN  553 => Ti := "100000010000001011100101111011111111000100010111"; --   -8322331   -1052393
      WHEN  554 => Ti := "100000010000111110101001111011111000110101100000"; --   -8319063   -1077920
      WHEN  555 => Ti := "100000010001110010111011111011110010100110110010"; --   -8315717   -1103438
      WHEN  556 => Ti := "100000010010101000011011111011101100011000001111"; --   -8312293   -1128945
      WHEN  557 => Ti := "100000010011011111001010111011100110001001110111"; --   -8308790   -1154441
      WHEN  558 => Ti := "100000010100010111000111111011011111111011101001"; --   -8305209   -1179927
      WHEN  559 => Ti := "100000010101010000010010111011011001101101100111"; --   -8301550   -1205401
      WHEN  560 => Ti := "100000010110001010101011111011010011011111110000"; --   -8297813   -1230864
      WHEN  561 => Ti := "100000010111000110010010111011001101010010000100"; --   -8293998   -1256316
      WHEN  562 => Ti := "100000011000000011001000111011000111000100100100"; --   -8290104   -1281756
      WHEN  563 => Ti := "100000011001000001001011111011000000110111010001"; --   -8286133   -1307183
      WHEN  564 => Ti := "100000011010000000011100111010111010101010001001"; --   -8282084   -1332599
      WHEN  565 => Ti := "100000011011000000111100111010110100011101001111"; --   -8277956   -1358001
      WHEN  566 => Ti := "100000011100000010101001111010101110010000100001"; --   -8273751   -1383391
      WHEN  567 => Ti := "100000011101000101100100111010101000000100000000"; --   -8269468   -1408768
      WHEN  568 => Ti := "100000011110001001101101111010100001110111101100"; --   -8265107   -1434132
      WHEN  569 => Ti := "100000011111001111000100111010011011101011100110"; --   -8260668   -1459482
      WHEN  570 => Ti := "100000100000010101101000111010010101011111101101"; --   -8256152   -1484819
      WHEN  571 => Ti := "100000100001011101011011111010001111010100000011"; --   -8251557   -1510141
      WHEN  572 => Ti := "100000100010100110011010111010001001001000100110"; --   -8246886   -1535450
      WHEN  573 => Ti := "100000100011110000101000111010000010111101011000"; --   -8242136   -1560744
      WHEN  574 => Ti := "100000100100111100000011111001111100110010011001"; --   -8237309   -1586023
      WHEN  575 => Ti := "100000100110001000101100111001110110100111101001"; --   -8232404   -1611287
      WHEN  576 => Ti := "100000100111010110100010111001110000011101001000"; --   -8227422   -1636536
      WHEN  577 => Ti := "100000101000100101100101111001101010010010110110"; --   -8222363   -1661770
      WHEN  578 => Ti := "100000101001110101110110111001100100001000110100"; --   -8217226   -1686988
      WHEN  579 => Ti := "100000101011000111010100111001011101111111000010"; --   -8212012   -1712190
      WHEN  580 => Ti := "100000101100011010000000111001010111110101100000"; --   -8206720   -1737376
      WHEN  581 => Ti := "100000101101101101111001111001010001101100001110"; --   -8201351   -1762546
      WHEN  582 => Ti := "100000101111000010111111111001001011100011001101"; --   -8195905   -1787699
      WHEN  583 => Ti := "100000110000011001010010111001000101011010011101"; --   -8190382   -1812835
      WHEN  584 => Ti := "100000110001110000110010111000111111010001111110"; --   -8184782   -1837954
      WHEN  585 => Ti := "100000110011001001100000111000111001001001110000"; --   -8179104   -1863056
      WHEN  586 => Ti := "100000110100100011011010111000110011000001110100"; --   -8173350   -1888140
      WHEN  587 => Ti := "100000110101111110100001111000101100111010001001"; --   -8167519   -1913207
      WHEN  588 => Ti := "100000110111011010110101111000100110110010110000"; --   -8161611   -1938256
      WHEN  589 => Ti := "100000111000111000010110111000100000101011101010"; --   -8155626   -1963286
      WHEN  590 => Ti := "100000111010010111000100111000011010100100110110"; --   -8149564   -1988298
      WHEN  591 => Ti := "100000111011110110111110111000010100011110010101"; --   -8143426   -2013291
      WHEN  592 => Ti := "100000111101011000000101111000001110011000000111"; --   -8137211   -2038265
      WHEN  593 => Ti := "100000111110111010011001111000001000010010001100"; --   -8130919   -2063220
      WHEN  594 => Ti := "100001000000011101111001111000000010001100100100"; --   -8124551   -2088156
      WHEN  595 => Ti := "100001000010000010100101110111111100000111010000"; --   -8118107   -2113072
      WHEN  596 => Ti := "100001000011101000011110110111110110000010010000"; --   -8111586   -2137968
      WHEN  597 => Ti := "100001000101001111100100110111101111111101100100"; --   -8104988   -2162844
      WHEN  598 => Ti := "100001000110110111110101110111101001111001001101"; --   -8098315   -2187699
      WHEN  599 => Ti := "100001001000100001010011110111100011110101001010"; --   -8091565   -2212534
      WHEN  600 => Ti := "100001001010001011111101110111011101110001011011"; --   -8084739   -2237349
      WHEN  601 => Ti := "100001001011110111110011110111010111101110000010"; --   -8077837   -2262142
      WHEN  602 => Ti := "100001001101100100110110110111010001101010111111"; --   -8070858   -2286913
      WHEN  603 => Ti := "100001001111010011000100110111001011101000010000"; --   -8063804   -2311664
      WHEN  604 => Ti := "100001010001000010011110110111000101100101111000"; --   -8056674   -2336392
      WHEN  605 => Ti := "100001010010110011000100110110111111100011110101"; --   -8049468   -2361099
      WHEN  606 => Ti := "100001010100100100110101110110111001100010001001"; --   -8042187   -2385783
      WHEN  607 => Ti := "100001010110010111110011110110110011100000110011"; --   -8034829   -2410445
      WHEN  608 => Ti := "100001011000001011111100110110101101011111110100"; --   -8027396   -2435084
      WHEN  609 => Ti := "100001011010000001010000110110100111011111001100"; --   -8019888   -2459700
      WHEN  610 => Ti := "100001011011110111110000110110100001011110111011"; --   -8012304   -2484293
      WHEN  611 => Ti := "100001011101101111011100110110011011011111000001"; --   -8004644   -2508863
      WHEN  612 => Ti := "100001011111101000010010110110010101011111011111"; --   -7996910   -2533409
      WHEN  613 => Ti := "100001100001100010010100110110001111100000010101"; --   -7989100   -2557931
      WHEN  614 => Ti := "100001100011011101100010110110001001100001100010"; --   -7981214   -2582430
      WHEN  615 => Ti := "100001100101011001111010110110000011100011001000"; --   -7973254   -2606904
      WHEN  616 => Ti := "100001100111010111011101110101111101100101000111"; --   -7965219   -2631353
      WHEN  617 => Ti := "100001101001010110001100110101110111100111011111"; --   -7957108   -2655777
      WHEN  618 => Ti := "100001101011010110000101110101110001101010001111"; --   -7948923   -2680177
      WHEN  619 => Ti := "100001101101010111001001110101101011101101011001"; --   -7940663   -2704551
      WHEN  620 => Ti := "100001101111011001011000110101100101110000111100"; --   -7932328   -2728900
      WHEN  621 => Ti := "100001110001011100110001110101011111110100111001"; --   -7923919   -2753223
      WHEN  622 => Ti := "100001110011100001010101110101011001111001001111"; --   -7915435   -2777521
      WHEN  623 => Ti := "100001110101100111000100110101010011111110000000"; --   -7906876   -2801792
      WHEN  624 => Ti := "100001110111101101111101110101001110000011001011"; --   -7898243   -2826037
      WHEN  625 => Ti := "100001111001110110000000110101001000001000110001"; --   -7889536   -2850255
      WHEN  626 => Ti := "100001111011111111001110110101000010001110110010"; --   -7880754   -2874446
      WHEN  627 => Ti := "100001111110001001100110110100111100010101001110"; --   -7871898   -2898610
      WHEN  628 => Ti := "100010000000010101000111110100110110011100000101"; --   -7862969   -2922747
      WHEN  629 => Ti := "100010000010100001110011110100110000100011010111"; --   -7853965   -2946857
      WHEN  630 => Ti := "100010000100101111101001110100101010101011000101"; --   -7844887   -2970939
      WHEN  631 => Ti := "100010000110111110101001110100100100110011010000"; --   -7835735   -2994992
      WHEN  632 => Ti := "100010001001001110110010110100011110111011110110"; --   -7826510   -3019018
      WHEN  633 => Ti := "100010001011100000000101110100011001000100111001"; --   -7817211   -3043015
      WHEN  634 => Ti := "100010001101110010100010110100010011001110011000"; --   -7807838   -3066984
      WHEN  635 => Ti := "100010010000000110001000110100001101011000010101"; --   -7798392   -3090923
      WHEN  636 => Ti := "100010010010011010110111110100000111100010101110"; --   -7788873   -3114834
      WHEN  637 => Ti := "100010010100110000110000110100000001101101100101"; --   -7779280   -3138715
      WHEN  638 => Ti := "100010010111000111110010110011111011111000111001"; --   -7769614   -3162567
      WHEN  639 => Ti := "100010011001011111111101110011110110000100101011"; --   -7759875   -3186389
      WHEN  640 => Ti := "100010011011111001010010110011110000010000111011"; --   -7750062   -3210181
      WHEN  641 => Ti := "100010011110010011101111110011101010011101101001"; --   -7740177   -3233943
      WHEN  642 => Ti := "100010100000101111010101110011100100101010110110"; --   -7730219   -3257674
      WHEN  643 => Ti := "100010100011001100000100110011011110111000100001"; --   -7720188   -3281375
      WHEN  644 => Ti := "100010100101101001111011110011011001000110101100"; --   -7710085   -3305044
      WHEN  645 => Ti := "100010101000001000111011110011010011010101010101"; --   -7699909   -3328683
      WHEN  646 => Ti := "100010101010101001000100110011001101100100011110"; --   -7689660   -3352290
      WHEN  647 => Ti := "100010101101001010010100110011000111110100000110"; --   -7679340   -3375866
      WHEN  648 => Ti := "100010101111101100101110110011000010000100001110"; --   -7668946   -3399410
      WHEN  649 => Ti := "100010110010010000001111110010111100010100110110"; --   -7658481   -3422922
      WHEN  650 => Ti := "100010110100110100111000110010110110100101111110"; --   -7647944   -3446402
      WHEN  651 => Ti := "100010110111011010101010110010110000110111100111"; --   -7637334   -3469849
      WHEN  652 => Ti := "100010111010000001100011110010101011001001110000"; --   -7626653   -3493264
      WHEN  653 => Ti := "100010111100101001100100110010100101011100011010"; --   -7615900   -3516646
      WHEN  654 => Ti := "100010111111010010101101110010011111101111100110"; --   -7605075   -3539994
      WHEN  655 => Ti := "100011000001111100111101110010011010000011010010"; --   -7594179   -3563310
      WHEN  656 => Ti := "100011000100101000010101110010010100010111100000"; --   -7583211   -3586592
      WHEN  657 => Ti := "100011000111010100110100110010001110101100010000"; --   -7572172   -3609840
      WHEN  658 => Ti := "100011001010000010011011110010001001000001100010"; --   -7561061   -3633054
      WHEN  659 => Ti := "100011001100110001001000110010000011010111010110"; --   -7549880   -3656234
      WHEN  660 => Ti := "100011001111100000111101110001111101101101101101"; --   -7538627   -3679379
      WHEN  661 => Ti := "100011010010010001111001110001111000000100100110"; --   -7527303   -3702490
      WHEN  662 => Ti := "100011010101000011111011110001110010011100000010"; --   -7515909   -3725566
      WHEN  663 => Ti := "100011010111110111000100110001101100110100000001"; --   -7504444   -3748607
      WHEN  664 => Ti := "100011011010101011010100110001100111001100100011"; --   -7492908   -3771613
      WHEN  665 => Ti := "100011011101100000101011110001100001100101101001"; --   -7481301   -3794583
      WHEN  666 => Ti := "100011100000010111001000110001011011111111010011"; --   -7469624   -3817517
      WHEN  667 => Ti := "100011100011001110101011110001010110011001100000"; --   -7457877   -3840416
      WHEN  668 => Ti := "100011100110000111010100110001010000110100010010"; --   -7446060   -3863278
      WHEN  669 => Ti := "100011101001000001000011110001001011001111101000"; --   -7434173   -3886104
      WHEN  670 => Ti := "100011101011111011111001110001000101101011100010"; --   -7422215   -3908894
      WHEN  671 => Ti := "100011101110110111110100110001000000001000000010"; --   -7410188   -3931646
      WHEN  672 => Ti := "100011110001110100110101110000111010100101000110"; --   -7398091   -3954362
      WHEN  673 => Ti := "100011110100110010111100110000110101000010110000"; --   -7385924   -3977040
      WHEN  674 => Ti := "100011110111110010001000110000101111100000111111"; --   -7373688   -3999681
      WHEN  675 => Ti := "100011111010110010011001110000101001111111110011"; --   -7361383   -4022285
      WHEN  676 => Ti := "100011111101110011110000110000100100011111001110"; --   -7349008   -4044850
      WHEN  677 => Ti := "100100000000110110001100110000011110111111001110"; --   -7336564   -4067378
      WHEN  678 => Ti := "100100000011111001101101110000011001011111110101"; --   -7324051   -4089867
      WHEN  679 => Ti := "100100000110111110010011110000010100000001000011"; --   -7311469   -4112317
      WHEN  680 => Ti := "100100001010000011111110110000001110100010110111"; --   -7298818   -4134729
      WHEN  681 => Ti := "100100001101001010101110110000001001000101010010"; --   -7286098   -4157102
      WHEN  682 => Ti := "100100010000010010100010110000000011101000010100"; --   -7273310   -4179436
      WHEN  683 => Ti := "100100010011011011011010101111111110001011111101"; --   -7260454   -4201731
      WHEN  684 => Ti := "100100010110100101010111101111111000110000001110"; --   -7247529   -4223986
      WHEN  685 => Ti := "100100011001110000011000101111110011010101000111"; --   -7234536   -4246201
      WHEN  686 => Ti := "100100011100111100011110101111101101111010101000"; --   -7221474   -4268376
      WHEN  687 => Ti := "100100100000001001100111101111101000100000110001"; --   -7208345   -4290511
      WHEN  688 => Ti := "100100100011010111110100101111100011000111100010"; --   -7195148   -4312606
      WHEN  689 => Ti := "100100100110100111000101101111011101101110111100"; --   -7181883   -4334660
      WHEN  690 => Ti := "100100101001110111011001101111011000010110111111"; --   -7168551   -4356673
      WHEN  691 => Ti := "100100101101001000110001101111010010111111101010"; --   -7155151   -4378646
      WHEN  692 => Ti := "100100110000011011001100101111001101101000111111"; --   -7141684   -4400577
      WHEN  693 => Ti := "100100110011101110101010101111001000010010111110"; --   -7128150   -4422466
      WHEN  694 => Ti := "100100110111000011001100101111000010111101100110"; --   -7114548   -4444314
      WHEN  695 => Ti := "100100111010011000110000101110111101101000110111"; --   -7100880   -4466121
      WHEN  696 => Ti := "100100111101101111010111101110111000010100110011"; --   -7087145   -4487885
      WHEN  697 => Ti := "100101000001000111000001101110110011000001011001"; --   -7073343   -4509607
      WHEN  698 => Ti := "100101000100011111101110101110101101101110101010"; --   -7059474   -4531286
      WHEN  699 => Ti := "100101000111111001011101101110101000011100100101"; --   -7045539   -4552923
      WHEN  700 => Ti := "100101001011010100001110101110100011001011001011"; --   -7031538   -4574517
      WHEN  701 => Ti := "100101001110110000000010101110011101111010011100"; --   -7017470   -4596068
      WHEN  702 => Ti := "100101010010001100110111101110011000101010011000"; --   -7003337   -4617576
      WHEN  703 => Ti := "100101010101101010101111101110010011011011000000"; --   -6989137   -4639040
      WHEN  704 => Ti := "100101011001001001101000101110001110001100010100"; --   -6974872   -4660460
      WHEN  705 => Ti := "100101011100101001100011101110001000111110010011"; --   -6960541   -4681837
      WHEN  706 => Ti := "100101100000001010100000101110000011110000111110"; --   -6946144   -4703170
      WHEN  707 => Ti := "100101100011101100011101101101111110100100010110"; --   -6931683   -4724458
      WHEN  708 => Ti := "100101100111001111011100101101111001011000011010"; --   -6917156   -4745702
      WHEN  709 => Ti := "100101101010110011011101101101110100001101001011"; --   -6902563   -4766901
      WHEN  710 => Ti := "100101101110011000011110101101101111000010101001"; --   -6887906   -4788055
      WHEN  711 => Ti := "100101110001111110100000101101101001111000110011"; --   -6873184   -4809165
      WHEN  712 => Ti := "100101110101100101100010101101100100101111101011"; --   -6858398   -4830229
      WHEN  713 => Ti := "100101111001001101100110101101011111100111010001"; --   -6843546   -4851247
      WHEN  714 => Ti := "100101111100110110101001101101011010011111100100"; --   -6828631   -4872220
      WHEN  715 => Ti := "100110000000100000101101101101010101011000100101"; --   -6813651   -4893147
      WHEN  716 => Ti := "100110000100001011110001101101010000010010010100"; --   -6798607   -4914028
      WHEN  717 => Ti := "100110000111110111110101101101001011001100110001"; --   -6783499   -4934863
      WHEN  718 => Ti := "100110001011100100111001101101000110000111111101"; --   -6768327   -4955651
      WHEN  719 => Ti := "100110001111010010111101101101000001000011110111"; --   -6753091   -4976393
      WHEN  720 => Ti := "100110010011000010000000101100111100000000100001"; --   -6737792   -4997087
      WHEN  721 => Ti := "100110010110110010000010101100110110111101111001"; --   -6722430   -5017735
      WHEN  722 => Ti := "100110011010100011000100101100110001111100000000"; --   -6707004   -5038336
      WHEN  723 => Ti := "100110011110010101000101101100101100111010110111"; --   -6691515   -5058889
      WHEN  724 => Ti := "100110100010001000000101101100100111111010011110"; --   -6675963   -5079394
      WHEN  725 => Ti := "100110100101111100000100101100100010111010110100"; --   -6660348   -5099852
      WHEN  726 => Ti := "100110101001110001000001101100011101111011111011"; --   -6644671   -5120261
      WHEN  727 => Ti := "100110101101100110111101101100011000111101110001"; --   -6628931   -5140623
      WHEN  728 => Ti := "100110110001011101111000101100010100000000011000"; --   -6613128   -5160936
      WHEN  729 => Ti := "100110110101010101110000101100001111000011101111"; --   -6597264   -5181201
      WHEN  730 => Ti := "100110111001001110100111101100001010000111111000"; --   -6581337   -5201416
      WHEN  731 => Ti := "100110111101001000011100101100000101001100110001"; --   -6565348   -5221583
      WHEN  732 => Ti := "100111000001000011001110101100000000010010011011"; --   -6549298   -5241701
      WHEN  733 => Ti := "100111000100111110111110101011111011011000110111"; --   -6533186   -5261769
      WHEN  734 => Ti := "100111001000111011101100101011110110100000000100"; --   -6517012   -5281788
      WHEN  735 => Ti := "100111001100111001010111101011110001101000000011"; --   -6500777   -5301757
      WHEN  736 => Ti := "100111010000110111111111101011101100110000110100"; --   -6484481   -5321676
      WHEN  737 => Ti := "100111010100110111100100101011100111111010010111"; --   -6468124   -5341545
      WHEN  738 => Ti := "100111011000111000000110101011100011000100101100"; --   -6451706   -5361364
      WHEN  739 => Ti := "100111011100111001100101101011011110001111110100"; --   -6435227   -5381132
      WHEN  740 => Ti := "100111100000111100000001101011011001011011101110"; --   -6418687   -5400850
      WHEN  741 => Ti := "100111100100111111011000101011010100101000011011"; --   -6402088   -5420517
      WHEN  742 => Ti := "100111101001000011101100101011001111110101111100"; --   -6385428   -5440132
      WHEN  743 => Ti := "100111101101001000111100101011001011000100001111"; --   -6368708   -5459697
      WHEN  744 => Ti := "100111110001001111001001101011000110010011010110"; --   -6351927   -5479210
      WHEN  745 => Ti := "100111110101010110010000101011000001100011010000"; --   -6335088   -5498672
      WHEN  746 => Ti := "100111111001011110010100101010111100110011111110"; --   -6318188   -5518082
      WHEN  747 => Ti := "100111111101100111010011101010111000000101100000"; --   -6301229   -5537440
      WHEN  748 => Ti := "101000000001110001001101101010110011010111110110"; --   -6284211   -5556746
      WHEN  749 => Ti := "101000000101111100000011101010101110101011000001"; --   -6267133   -5575999
      WHEN  750 => Ti := "101000001010000111110011101010101001111111000000"; --   -6249997   -5595200
      WHEN  751 => Ti := "101000001110010100011110101010100101010011110011"; --   -6232802   -5614349
      WHEN  752 => Ti := "101000010010100010000100101010100000101001011100"; --   -6215548   -5633444
      WHEN  753 => Ti := "101000010110110000100101101010011011111111111001"; --   -6198235   -5652487
      WHEN  754 => Ti := "101000011010111111111111101010010111010111001100"; --   -6180865   -5671476
      WHEN  755 => Ti := "101000011111010000010100101010010010101111010100"; --   -6163436   -5690412
      WHEN  756 => Ti := "101000100011100001100011101010001110001000010010"; --   -6145949   -5709294
      WHEN  757 => Ti := "101000100111110011101100101010001001100010000101"; --   -6128404   -5728123
      WHEN  758 => Ti := "101000101100000110101111101010000100111100101110"; --   -6110801   -5746898
      WHEN  759 => Ti := "101000110000011010101011101010000000011000001110"; --   -6093141   -5765618
      WHEN  760 => Ti := "101000110100101111100000101001111011110100100011"; --   -6075424   -5784285
      WHEN  761 => Ti := "101000111001000101001110101001110111010001101111"; --   -6057650   -5802897
      WHEN  762 => Ti := "101000111101011011110110101001110010101111110010"; --   -6039818   -5821454
      WHEN  763 => Ti := "101001000001110011010110101001101110001110101100"; --   -6021930   -5839956
      WHEN  764 => Ti := "101001000110001011101111101001101001101110011100"; --   -6003985   -5858404
      WHEN  765 => Ti := "101001001010100101000001101001100101001111000100"; --   -5985983   -5876796
      WHEN  766 => Ti := "101001001110111111001011101001100000110000100011"; --   -5967925   -5895133
      WHEN  767 => Ti := "101001010011011010001101101001011100010010111001"; --   -5949811   -5913415
      WHEN  768 => Ti := "101001010111110110000111101001010111110110000111"; --   -5931641   -5931641
      WHEN  769 => Ti := "101001011100010010111001101001010011011010001101"; --   -5913415   -5949811
      WHEN  770 => Ti := "101001100000110000100011101001001110111111001011"; --   -5895133   -5967925
      WHEN  771 => Ti := "101001100101001111000100101001001010100101000001"; --   -5876796   -5985983
      WHEN  772 => Ti := "101001101001101110011100101001000110001011101111"; --   -5858404   -6003985
      WHEN  773 => Ti := "101001101110001110101100101001000001110011010110"; --   -5839956   -6021930
      WHEN  774 => Ti := "101001110010101111110010101000111101011011110110"; --   -5821454   -6039818
      WHEN  775 => Ti := "101001110111010001101111101000111001000101001110"; --   -5802897   -6057650
      WHEN  776 => Ti := "101001111011110100100011101000110100101111100000"; --   -5784285   -6075424
      WHEN  777 => Ti := "101010000000011000001110101000110000011010101011"; --   -5765618   -6093141
      WHEN  778 => Ti := "101010000100111100101110101000101100000110101111"; --   -5746898   -6110801
      WHEN  779 => Ti := "101010001001100010000101101000100111110011101100"; --   -5728123   -6128404
      WHEN  780 => Ti := "101010001110001000010010101000100011100001100011"; --   -5709294   -6145949
      WHEN  781 => Ti := "101010010010101111010100101000011111010000010100"; --   -5690412   -6163436
      WHEN  782 => Ti := "101010010111010111001100101000011010111111111111"; --   -5671476   -6180865
      WHEN  783 => Ti := "101010011011111111111001101000010110110000100101"; --   -5652487   -6198235
      WHEN  784 => Ti := "101010100000101001011100101000010010100010000100"; --   -5633444   -6215548
      WHEN  785 => Ti := "101010100101010011110011101000001110010100011110"; --   -5614349   -6232802
      WHEN  786 => Ti := "101010101001111111000000101000001010000111110011"; --   -5595200   -6249997
      WHEN  787 => Ti := "101010101110101011000001101000000101111100000011"; --   -5575999   -6267133
      WHEN  788 => Ti := "101010110011010111110110101000000001110001001101"; --   -5556746   -6284211
      WHEN  789 => Ti := "101010111000000101100000100111111101100111010011"; --   -5537440   -6301229
      WHEN  790 => Ti := "101010111100110011111110100111111001011110010100"; --   -5518082   -6318188
      WHEN  791 => Ti := "101011000001100011010000100111110101010110010000"; --   -5498672   -6335088
      WHEN  792 => Ti := "101011000110010011010110100111110001001111001001"; --   -5479210   -6351927
      WHEN  793 => Ti := "101011001011000100001111100111101101001000111100"; --   -5459697   -6368708
      WHEN  794 => Ti := "101011001111110101111100100111101001000011101100"; --   -5440132   -6385428
      WHEN  795 => Ti := "101011010100101000011011100111100100111111011000"; --   -5420517   -6402088
      WHEN  796 => Ti := "101011011001011011101110100111100000111100000001"; --   -5400850   -6418687
      WHEN  797 => Ti := "101011011110001111110100100111011100111001100101"; --   -5381132   -6435227
      WHEN  798 => Ti := "101011100011000100101100100111011000111000000110"; --   -5361364   -6451706
      WHEN  799 => Ti := "101011100111111010010111100111010100110111100100"; --   -5341545   -6468124
      WHEN  800 => Ti := "101011101100110000110100100111010000110111111111"; --   -5321676   -6484481
      WHEN  801 => Ti := "101011110001101000000011100111001100111001010111"; --   -5301757   -6500777
      WHEN  802 => Ti := "101011110110100000000100100111001000111011101100"; --   -5281788   -6517012
      WHEN  803 => Ti := "101011111011011000110111100111000100111110111110"; --   -5261769   -6533186
      WHEN  804 => Ti := "101100000000010010011011100111000001000011001110"; --   -5241701   -6549298
      WHEN  805 => Ti := "101100000101001100110001100110111101001000011100"; --   -5221583   -6565348
      WHEN  806 => Ti := "101100001010000111111000100110111001001110100111"; --   -5201416   -6581337
      WHEN  807 => Ti := "101100001111000011101111100110110101010101110000"; --   -5181201   -6597264
      WHEN  808 => Ti := "101100010100000000011000100110110001011101111000"; --   -5160936   -6613128
      WHEN  809 => Ti := "101100011000111101110001100110101101100110111101"; --   -5140623   -6628931
      WHEN  810 => Ti := "101100011101111011111011100110101001110001000001"; --   -5120261   -6644671
      WHEN  811 => Ti := "101100100010111010110100100110100101111100000100"; --   -5099852   -6660348
      WHEN  812 => Ti := "101100100111111010011110100110100010001000000101"; --   -5079394   -6675963
      WHEN  813 => Ti := "101100101100111010110111100110011110010101000101"; --   -5058889   -6691515
      WHEN  814 => Ti := "101100110001111100000000100110011010100011000100"; --   -5038336   -6707004
      WHEN  815 => Ti := "101100110110111101111001100110010110110010000010"; --   -5017735   -6722430
      WHEN  816 => Ti := "101100111100000000100001100110010011000010000000"; --   -4997087   -6737792
      WHEN  817 => Ti := "101101000001000011110111100110001111010010111101"; --   -4976393   -6753091
      WHEN  818 => Ti := "101101000110000111111101100110001011100100111001"; --   -4955651   -6768327
      WHEN  819 => Ti := "101101001011001100110001100110000111110111110101"; --   -4934863   -6783499
      WHEN  820 => Ti := "101101010000010010010100100110000100001011110001"; --   -4914028   -6798607
      WHEN  821 => Ti := "101101010101011000100101100110000000100000101101"; --   -4893147   -6813651
      WHEN  822 => Ti := "101101011010011111100100100101111100110110101001"; --   -4872220   -6828631
      WHEN  823 => Ti := "101101011111100111010001100101111001001101100110"; --   -4851247   -6843546
      WHEN  824 => Ti := "101101100100101111101011100101110101100101100010"; --   -4830229   -6858398
      WHEN  825 => Ti := "101101101001111000110011100101110001111110100000"; --   -4809165   -6873184
      WHEN  826 => Ti := "101101101111000010101001100101101110011000011110"; --   -4788055   -6887906
      WHEN  827 => Ti := "101101110100001101001011100101101010110011011101"; --   -4766901   -6902563
      WHEN  828 => Ti := "101101111001011000011010100101100111001111011100"; --   -4745702   -6917156
      WHEN  829 => Ti := "101101111110100100010110100101100011101100011101"; --   -4724458   -6931683
      WHEN  830 => Ti := "101110000011110000111110100101100000001010100000"; --   -4703170   -6946144
      WHEN  831 => Ti := "101110001000111110010011100101011100101001100011"; --   -4681837   -6960541
      WHEN  832 => Ti := "101110001110001100010100100101011001001001101000"; --   -4660460   -6974872
      WHEN  833 => Ti := "101110010011011011000000100101010101101010101111"; --   -4639040   -6989137
      WHEN  834 => Ti := "101110011000101010011000100101010010001100110111"; --   -4617576   -7003337
      WHEN  835 => Ti := "101110011101111010011100100101001110110000000010"; --   -4596068   -7017470
      WHEN  836 => Ti := "101110100011001011001011100101001011010100001110"; --   -4574517   -7031538
      WHEN  837 => Ti := "101110101000011100100101100101000111111001011101"; --   -4552923   -7045539
      WHEN  838 => Ti := "101110101101101110101010100101000100011111101110"; --   -4531286   -7059474
      WHEN  839 => Ti := "101110110011000001011001100101000001000111000001"; --   -4509607   -7073343
      WHEN  840 => Ti := "101110111000010100110011100100111101101111010111"; --   -4487885   -7087145
      WHEN  841 => Ti := "101110111101101000110111100100111010011000110000"; --   -4466121   -7100880
      WHEN  842 => Ti := "101111000010111101100110100100110111000011001100"; --   -4444314   -7114548
      WHEN  843 => Ti := "101111001000010010111110100100110011101110101010"; --   -4422466   -7128150
      WHEN  844 => Ti := "101111001101101000111111100100110000011011001100"; --   -4400577   -7141684
      WHEN  845 => Ti := "101111010010111111101010100100101101001000110001"; --   -4378646   -7155151
      WHEN  846 => Ti := "101111011000010110111111100100101001110111011001"; --   -4356673   -7168551
      WHEN  847 => Ti := "101111011101101110111100100100100110100111000101"; --   -4334660   -7181883
      WHEN  848 => Ti := "101111100011000111100010100100100011010111110100"; --   -4312606   -7195148
      WHEN  849 => Ti := "101111101000100000110001100100100000001001100111"; --   -4290511   -7208345
      WHEN  850 => Ti := "101111101101111010101000100100011100111100011110"; --   -4268376   -7221474
      WHEN  851 => Ti := "101111110011010101000111100100011001110000011000"; --   -4246201   -7234536
      WHEN  852 => Ti := "101111111000110000001110100100010110100101010111"; --   -4223986   -7247529
      WHEN  853 => Ti := "101111111110001011111101100100010011011011011010"; --   -4201731   -7260454
      WHEN  854 => Ti := "110000000011101000010100100100010000010010100010"; --   -4179436   -7273310
      WHEN  855 => Ti := "110000001001000101010010100100001101001010101110"; --   -4157102   -7286098
      WHEN  856 => Ti := "110000001110100010110111100100001010000011111110"; --   -4134729   -7298818
      WHEN  857 => Ti := "110000010100000001000011100100000110111110010011"; --   -4112317   -7311469
      WHEN  858 => Ti := "110000011001011111110101100100000011111001101101"; --   -4089867   -7324051
      WHEN  859 => Ti := "110000011110111111001110100100000000110110001100"; --   -4067378   -7336564
      WHEN  860 => Ti := "110000100100011111001110100011111101110011110000"; --   -4044850   -7349008
      WHEN  861 => Ti := "110000101001111111110011100011111010110010011001"; --   -4022285   -7361383
      WHEN  862 => Ti := "110000101111100000111111100011110111110010001000"; --   -3999681   -7373688
      WHEN  863 => Ti := "110000110101000010110000100011110100110010111100"; --   -3977040   -7385924
      WHEN  864 => Ti := "110000111010100101000110100011110001110100110101"; --   -3954362   -7398091
      WHEN  865 => Ti := "110001000000001000000010100011101110110111110100"; --   -3931646   -7410188
      WHEN  866 => Ti := "110001000101101011100010100011101011111011111001"; --   -3908894   -7422215
      WHEN  867 => Ti := "110001001011001111101000100011101001000001000011"; --   -3886104   -7434173
      WHEN  868 => Ti := "110001010000110100010010100011100110000111010100"; --   -3863278   -7446060
      WHEN  869 => Ti := "110001010110011001100000100011100011001110101011"; --   -3840416   -7457877
      WHEN  870 => Ti := "110001011011111111010011100011100000010111001000"; --   -3817517   -7469624
      WHEN  871 => Ti := "110001100001100101101001100011011101100000101011"; --   -3794583   -7481301
      WHEN  872 => Ti := "110001100111001100100011100011011010101011010100"; --   -3771613   -7492908
      WHEN  873 => Ti := "110001101100110100000001100011010111110111000100"; --   -3748607   -7504444
      WHEN  874 => Ti := "110001110010011100000010100011010101000011111011"; --   -3725566   -7515909
      WHEN  875 => Ti := "110001111000000100100110100011010010010001111001"; --   -3702490   -7527303
      WHEN  876 => Ti := "110001111101101101101101100011001111100000111101"; --   -3679379   -7538627
      WHEN  877 => Ti := "110010000011010111010110100011001100110001001000"; --   -3656234   -7549880
      WHEN  878 => Ti := "110010001001000001100010100011001010000010011011"; --   -3633054   -7561061
      WHEN  879 => Ti := "110010001110101100010000100011000111010100110100"; --   -3609840   -7572172
      WHEN  880 => Ti := "110010010100010111100000100011000100101000010101"; --   -3586592   -7583211
      WHEN  881 => Ti := "110010011010000011010010100011000001111100111101"; --   -3563310   -7594179
      WHEN  882 => Ti := "110010011111101111100110100010111111010010101101"; --   -3539994   -7605075
      WHEN  883 => Ti := "110010100101011100011010100010111100101001100100"; --   -3516646   -7615900
      WHEN  884 => Ti := "110010101011001001110000100010111010000001100011"; --   -3493264   -7626653
      WHEN  885 => Ti := "110010110000110111100111100010110111011010101010"; --   -3469849   -7637334
      WHEN  886 => Ti := "110010110110100101111110100010110100110100111000"; --   -3446402   -7647944
      WHEN  887 => Ti := "110010111100010100110110100010110010010000001111"; --   -3422922   -7658481
      WHEN  888 => Ti := "110011000010000100001110100010101111101100101110"; --   -3399410   -7668946
      WHEN  889 => Ti := "110011000111110100000110100010101101001010010100"; --   -3375866   -7679340
      WHEN  890 => Ti := "110011001101100100011110100010101010101001000100"; --   -3352290   -7689660
      WHEN  891 => Ti := "110011010011010101010101100010101000001000111011"; --   -3328683   -7699909
      WHEN  892 => Ti := "110011011001000110101100100010100101101001111011"; --   -3305044   -7710085
      WHEN  893 => Ti := "110011011110111000100001100010100011001100000100"; --   -3281375   -7720188
      WHEN  894 => Ti := "110011100100101010110110100010100000101111010101"; --   -3257674   -7730219
      WHEN  895 => Ti := "110011101010011101101001100010011110010011101111"; --   -3233943   -7740177
      WHEN  896 => Ti := "110011110000010000111011100010011011111001010010"; --   -3210181   -7750062
      WHEN  897 => Ti := "110011110110000100101011100010011001011111111101"; --   -3186389   -7759875
      WHEN  898 => Ti := "110011111011111000111001100010010111000111110010"; --   -3162567   -7769614
      WHEN  899 => Ti := "110100000001101101100101100010010100110000110000"; --   -3138715   -7779280
      WHEN  900 => Ti := "110100000111100010101110100010010010011010110111"; --   -3114834   -7788873
      WHEN  901 => Ti := "110100001101011000010101100010010000000110001000"; --   -3090923   -7798392
      WHEN  902 => Ti := "110100010011001110011000100010001101110010100010"; --   -3066984   -7807838
      WHEN  903 => Ti := "110100011001000100111001100010001011100000000101"; --   -3043015   -7817211
      WHEN  904 => Ti := "110100011110111011110110100010001001001110110010"; --   -3019018   -7826510
      WHEN  905 => Ti := "110100100100110011010000100010000110111110101001"; --   -2994992   -7835735
      WHEN  906 => Ti := "110100101010101011000101100010000100101111101001"; --   -2970939   -7844887
      WHEN  907 => Ti := "110100110000100011010111100010000010100001110011"; --   -2946857   -7853965
      WHEN  908 => Ti := "110100110110011100000101100010000000010101000111"; --   -2922747   -7862969
      WHEN  909 => Ti := "110100111100010101001110100001111110001001100110"; --   -2898610   -7871898
      WHEN  910 => Ti := "110101000010001110110010100001111011111111001110"; --   -2874446   -7880754
      WHEN  911 => Ti := "110101001000001000110001100001111001110110000000"; --   -2850255   -7889536
      WHEN  912 => Ti := "110101001110000011001011100001110111101101111101"; --   -2826037   -7898243
      WHEN  913 => Ti := "110101010011111110000000100001110101100111000100"; --   -2801792   -7906876
      WHEN  914 => Ti := "110101011001111001001111100001110011100001010101"; --   -2777521   -7915435
      WHEN  915 => Ti := "110101011111110100111001100001110001011100110001"; --   -2753223   -7923919
      WHEN  916 => Ti := "110101100101110000111100100001101111011001011000"; --   -2728900   -7932328
      WHEN  917 => Ti := "110101101011101101011001100001101101010111001001"; --   -2704551   -7940663
      WHEN  918 => Ti := "110101110001101010001111100001101011010110000101"; --   -2680177   -7948923
      WHEN  919 => Ti := "110101110111100111011111100001101001010110001100"; --   -2655777   -7957108
      WHEN  920 => Ti := "110101111101100101000111100001100111010111011101"; --   -2631353   -7965219
      WHEN  921 => Ti := "110110000011100011001000100001100101011001111010"; --   -2606904   -7973254
      WHEN  922 => Ti := "110110001001100001100010100001100011011101100010"; --   -2582430   -7981214
      WHEN  923 => Ti := "110110001111100000010101100001100001100010010100"; --   -2557931   -7989100
      WHEN  924 => Ti := "110110010101011111011111100001011111101000010010"; --   -2533409   -7996910
      WHEN  925 => Ti := "110110011011011111000001100001011101101111011100"; --   -2508863   -8004644
      WHEN  926 => Ti := "110110100001011110111011100001011011110111110000"; --   -2484293   -8012304
      WHEN  927 => Ti := "110110100111011111001100100001011010000001010000"; --   -2459700   -8019888
      WHEN  928 => Ti := "110110101101011111110100100001011000001011111100"; --   -2435084   -8027396
      WHEN  929 => Ti := "110110110011100000110011100001010110010111110011"; --   -2410445   -8034829
      WHEN  930 => Ti := "110110111001100010001001100001010100100100110101"; --   -2385783   -8042187
      WHEN  931 => Ti := "110110111111100011110101100001010010110011000100"; --   -2361099   -8049468
      WHEN  932 => Ti := "110111000101100101111000100001010001000010011110"; --   -2336392   -8056674
      WHEN  933 => Ti := "110111001011101000010000100001001111010011000100"; --   -2311664   -8063804
      WHEN  934 => Ti := "110111010001101010111111100001001101100100110110"; --   -2286913   -8070858
      WHEN  935 => Ti := "110111010111101110000010100001001011110111110011"; --   -2262142   -8077837
      WHEN  936 => Ti := "110111011101110001011011100001001010001011111101"; --   -2237349   -8084739
      WHEN  937 => Ti := "110111100011110101001010100001001000100001010011"; --   -2212534   -8091565
      WHEN  938 => Ti := "110111101001111001001101100001000110110111110101"; --   -2187699   -8098315
      WHEN  939 => Ti := "110111101111111101100100100001000101001111100100"; --   -2162844   -8104988
      WHEN  940 => Ti := "110111110110000010010000100001000011101000011110"; --   -2137968   -8111586
      WHEN  941 => Ti := "110111111100000111010000100001000010000010100101"; --   -2113072   -8118107
      WHEN  942 => Ti := "111000000010001100100100100001000000011101111001"; --   -2088156   -8124551
      WHEN  943 => Ti := "111000001000010010001100100000111110111010011001"; --   -2063220   -8130919
      WHEN  944 => Ti := "111000001110011000000111100000111101011000000101"; --   -2038265   -8137211
      WHEN  945 => Ti := "111000010100011110010101100000111011110110111110"; --   -2013291   -8143426
      WHEN  946 => Ti := "111000011010100100110110100000111010010111000100"; --   -1988298   -8149564
      WHEN  947 => Ti := "111000100000101011101010100000111000111000010110"; --   -1963286   -8155626
      WHEN  948 => Ti := "111000100110110010110000100000110111011010110101"; --   -1938256   -8161611
      WHEN  949 => Ti := "111000101100111010001001100000110101111110100001"; --   -1913207   -8167519
      WHEN  950 => Ti := "111000110011000001110100100000110100100011011010"; --   -1888140   -8173350
      WHEN  951 => Ti := "111000111001001001110000100000110011001001100000"; --   -1863056   -8179104
      WHEN  952 => Ti := "111000111111010001111110100000110001110000110010"; --   -1837954   -8184782
      WHEN  953 => Ti := "111001000101011010011101100000110000011001010010"; --   -1812835   -8190382
      WHEN  954 => Ti := "111001001011100011001101100000101111000010111111"; --   -1787699   -8195905
      WHEN  955 => Ti := "111001010001101100001110100000101101101101111001"; --   -1762546   -8201351
      WHEN  956 => Ti := "111001010111110101100000100000101100011010000000"; --   -1737376   -8206720
      WHEN  957 => Ti := "111001011101111111000010100000101011000111010100"; --   -1712190   -8212012
      WHEN  958 => Ti := "111001100100001000110100100000101001110101110110"; --   -1686988   -8217226
      WHEN  959 => Ti := "111001101010010010110110100000101000100101100101"; --   -1661770   -8222363
      WHEN  960 => Ti := "111001110000011101001000100000100111010110100010"; --   -1636536   -8227422
      WHEN  961 => Ti := "111001110110100111101001100000100110001000101100"; --   -1611287   -8232404
      WHEN  962 => Ti := "111001111100110010011001100000100100111100000011"; --   -1586023   -8237309
      WHEN  963 => Ti := "111010000010111101011000100000100011110000101000"; --   -1560744   -8242136
      WHEN  964 => Ti := "111010001001001000100110100000100010100110011010"; --   -1535450   -8246886
      WHEN  965 => Ti := "111010001111010100000011100000100001011101011011"; --   -1510141   -8251557
      WHEN  966 => Ti := "111010010101011111101101100000100000010101101000"; --   -1484819   -8256152
      WHEN  967 => Ti := "111010011011101011100110100000011111001111000100"; --   -1459482   -8260668
      WHEN  968 => Ti := "111010100001110111101100100000011110001001101101"; --   -1434132   -8265107
      WHEN  969 => Ti := "111010101000000100000000100000011101000101100100"; --   -1408768   -8269468
      WHEN  970 => Ti := "111010101110010000100001100000011100000010101001"; --   -1383391   -8273751
      WHEN  971 => Ti := "111010110100011101001111100000011011000000111100"; --   -1358001   -8277956
      WHEN  972 => Ti := "111010111010101010001001100000011010000000011100"; --   -1332599   -8282084
      WHEN  973 => Ti := "111011000000110111010001100000011001000001001011"; --   -1307183   -8286133
      WHEN  974 => Ti := "111011000111000100100100100000011000000011001000"; --   -1281756   -8290104
      WHEN  975 => Ti := "111011001101010010000100100000010111000110010010"; --   -1256316   -8293998
      WHEN  976 => Ti := "111011010011011111110000100000010110001010101011"; --   -1230864   -8297813
      WHEN  977 => Ti := "111011011001101101100111100000010101010000010010"; --   -1205401   -8301550
      WHEN  978 => Ti := "111011011111111011101001100000010100010111000111"; --   -1179927   -8305209
      WHEN  979 => Ti := "111011100110001001110111100000010011011111001010"; --   -1154441   -8308790
      WHEN  980 => Ti := "111011101100011000001111100000010010101000011011"; --   -1128945   -8312293
      WHEN  981 => Ti := "111011110010100110110010100000010001110010111011"; --   -1103438   -8315717
      WHEN  982 => Ti := "111011111000110101100000100000010000111110101001"; --   -1077920   -8319063
      WHEN  983 => Ti := "111011111111000100010111100000010000001011100101"; --   -1052393   -8322331
      WHEN  984 => Ti := "111100000101010011011001100000001111011001101111"; --   -1026855   -8325521
      WHEN  985 => Ti := "111100001011100010100100100000001110101001001000"; --   -1001308   -8328632
      WHEN  986 => Ti := "111100010001110001111001100000001101111001101111"; --    -975751   -8331665
      WHEN  987 => Ti := "111100011000000001010110100000001101001011100101"; --    -950186   -8334619
      WHEN  988 => Ti := "111100011110010000111101100000001100011110101001"; --    -924611   -8337495
      WHEN  989 => Ti := "111100100100100000101101100000001011110010111100"; --    -899027   -8340292
      WHEN  990 => Ti := "111100101010110000100101100000001011001000011101"; --    -873435   -8343011
      WHEN  991 => Ti := "111100110001000000100101100000001010011111001100"; --    -847835   -8345652
      WHEN  992 => Ti := "111100110111010000101101100000001001110111001010"; --    -822227   -8348214
      WHEN  993 => Ti := "111100111101100000111101100000001001010000010111"; --    -796611   -8350697
      WHEN  994 => Ti := "111101000011110001010100100000001000101010110010"; --    -770988   -8353102
      WHEN  995 => Ti := "111101001010000001110010100000001000000110011100"; --    -745358   -8355428
      WHEN  996 => Ti := "111101010000010010011000100000000111100011010101"; --    -719720   -8357675
      WHEN  997 => Ti := "111101010110100011000100100000000111000001011100"; --    -694076   -8359844
      WHEN  998 => Ti := "111101011100110011110111100000000110100000110010"; --    -668425   -8361934
      WHEN  999 => Ti := "111101100011000100110001100000000110000001010111"; --    -642767   -8363945
      WHEN 1000 => Ti := "111101101001010101110000100000000101100011001010"; --    -617104   -8365878
      WHEN 1001 => Ti := "111101101111100110110101100000000101000110001100"; --    -591435   -8367732
      WHEN 1002 => Ti := "111101110101110111111111100000000100101010011101"; --    -565761   -8369507
      WHEN 1003 => Ti := "111101111100001001001111100000000100001111111101"; --    -540081   -8371203
      WHEN 1004 => Ti := "111110000010011010100100100000000011110110101011"; --    -514396   -8372821
      WHEN 1005 => Ti := "111110001000101011111110100000000011011110101001"; --    -488706   -8374359
      WHEN 1006 => Ti := "111110001110111101011101100000000011000111110101"; --    -463011   -8375819
      WHEN 1007 => Ti := "111110010101001111000000100000000010110010010000"; --    -437312   -8377200
      WHEN 1008 => Ti := "111110011011100000100111100000000010011101111001"; --    -411609   -8378503
      WHEN 1009 => Ti := "111110100001110010010001100000000010001010110010"; --    -385903   -8379726
      WHEN 1010 => Ti := "111110101000000100000000100000000001111000111010"; --    -360192   -8380870
      WHEN 1011 => Ti := "111110101110010101110010100000000001101000010000"; --    -334478   -8381936
      WHEN 1012 => Ti := "111110110100100111100111100000000001011000110101"; --    -308761   -8382923
      WHEN 1013 => Ti := "111110111010111001011111100000000001001010101001"; --    -283041   -8383831
      WHEN 1014 => Ti := "111111000001001011011001100000000000111101101101"; --    -257319   -8384659
      WHEN 1015 => Ti := "111111000111011101010110100000000000110001111111"; --    -231594   -8385409
      WHEN 1016 => Ti := "111111001101101111010101100000000000100111011111"; --    -205867   -8386081
      WHEN 1017 => Ti := "111111010100000001010110100000000000011110001111"; --    -180138   -8386673
      WHEN 1018 => Ti := "111111011010010011011001100000000000010110001110"; --    -154407   -8387186
      WHEN 1019 => Ti := "111111100000100101011101100000000000001111011100"; --    -128675   -8387620
      WHEN 1020 => Ti := "111111100110110111100011100000000000001001111001"; --    -102941   -8387975
      WHEN 1021 => Ti := "111111101101001001101001100000000000000101100100"; --     -77207   -8388252
      WHEN 1022 => Ti := "111111110011011011110000100000000000000010011111"; --     -51472   -8388449
      WHEN 1023 => Ti := "111111111001101101111000100000000000000000101000"; --     -25736   -8388568
      WHEN OTHERS => Ti := "000000000000000000000000011111111111111111111111"; --         +0   +8388607
    END CASE; 
    T <= Ti; 
  END PROCESS; 
END ARCHITECTURE rtl; 
